magic
tech scmos
timestamp 1684763702
<< ab >>
rect -547 6 -467 77
rect -464 6 -424 77
rect -360 6 -320 77
rect -318 6 -278 77
rect -274 6 -234 77
rect -205 6 -165 77
rect -161 6 -121 77
rect -119 6 -79 77
rect -78 6 -38 77
rect -35 6 45 77
rect 48 6 88 77
rect -582 5 -395 6
rect -582 -66 -486 5
rect -483 -66 -395 5
rect -394 5 88 6
rect -394 -66 -266 5
rect -265 -66 -177 5
rect -176 -66 -48 5
rect -44 -66 52 5
rect -519 -138 -431 -66
rect -430 -138 -302 -66
rect -299 -138 -211 -66
rect -210 -138 11 -66
<< nwell >>
rect -552 37 93 82
rect -587 -71 57 -26
rect -524 -106 16 -71
<< pwell >>
rect -552 11 93 37
rect -587 0 93 11
rect -587 -26 57 0
rect -524 -143 16 -106
<< poly >>
rect -538 62 -536 66
rect -528 64 -526 69
rect -518 64 -516 69
rect -498 62 -496 66
rect -488 64 -486 69
rect -478 64 -476 69
rect -538 40 -536 44
rect -528 40 -526 51
rect -518 48 -516 51
rect -518 46 -512 48
rect -518 44 -516 46
rect -514 44 -512 46
rect -455 62 -453 66
rect -445 64 -443 69
rect -435 64 -433 69
rect -518 42 -512 44
rect -538 38 -532 40
rect -538 36 -536 38
rect -534 36 -532 38
rect -538 34 -532 36
rect -528 38 -522 40
rect -528 36 -526 38
rect -524 36 -522 38
rect -528 34 -522 36
rect -538 29 -536 34
rect -525 29 -523 34
rect -518 29 -516 42
rect -498 40 -496 44
rect -488 40 -486 51
rect -478 48 -476 51
rect -478 46 -472 48
rect -478 44 -476 46
rect -474 44 -472 46
rect -351 62 -349 66
rect -341 64 -339 69
rect -331 64 -329 69
rect -478 42 -472 44
rect -498 38 -492 40
rect -498 36 -496 38
rect -494 36 -492 38
rect -498 34 -492 36
rect -488 38 -482 40
rect -488 36 -486 38
rect -484 36 -482 38
rect -488 34 -482 36
rect -498 29 -496 34
rect -485 29 -483 34
rect -478 29 -476 42
rect -455 40 -453 44
rect -445 40 -443 51
rect -435 48 -433 51
rect -435 46 -429 48
rect -435 44 -433 46
rect -431 44 -429 46
rect -309 62 -307 66
rect -299 64 -297 69
rect -289 64 -287 69
rect -435 42 -429 44
rect -455 38 -449 40
rect -455 36 -453 38
rect -451 36 -449 38
rect -455 34 -449 36
rect -445 38 -439 40
rect -445 36 -443 38
rect -441 36 -439 38
rect -445 34 -439 36
rect -455 29 -453 34
rect -442 29 -440 34
rect -435 29 -433 42
rect -351 40 -349 44
rect -341 40 -339 51
rect -331 48 -329 51
rect -331 46 -325 48
rect -331 44 -329 46
rect -327 44 -325 46
rect -265 62 -263 66
rect -255 64 -253 69
rect -245 64 -243 69
rect -331 42 -325 44
rect -351 38 -345 40
rect -351 36 -349 38
rect -347 36 -345 38
rect -351 34 -345 36
rect -341 38 -335 40
rect -341 36 -339 38
rect -337 36 -335 38
rect -341 34 -335 36
rect -351 29 -349 34
rect -338 29 -336 34
rect -331 29 -329 42
rect -309 40 -307 44
rect -299 40 -297 51
rect -289 48 -287 51
rect -289 46 -283 48
rect -289 44 -287 46
rect -285 44 -283 46
rect -196 62 -194 66
rect -186 64 -184 69
rect -176 64 -174 69
rect -289 42 -283 44
rect -309 38 -303 40
rect -309 36 -307 38
rect -305 36 -303 38
rect -309 34 -303 36
rect -299 38 -293 40
rect -299 36 -297 38
rect -295 36 -293 38
rect -299 34 -293 36
rect -309 29 -307 34
rect -296 29 -294 34
rect -289 29 -287 42
rect -265 40 -263 44
rect -255 40 -253 51
rect -245 48 -243 51
rect -245 46 -239 48
rect -245 44 -243 46
rect -241 44 -239 46
rect -152 62 -150 66
rect -142 64 -140 69
rect -132 64 -130 69
rect -245 42 -239 44
rect -265 38 -259 40
rect -265 36 -263 38
rect -261 36 -259 38
rect -265 34 -259 36
rect -255 38 -249 40
rect -255 36 -253 38
rect -251 36 -249 38
rect -255 34 -249 36
rect -265 29 -263 34
rect -252 29 -250 34
rect -245 29 -243 42
rect -196 40 -194 44
rect -186 40 -184 51
rect -176 48 -174 51
rect -176 46 -170 48
rect -176 44 -174 46
rect -172 44 -170 46
rect -110 62 -108 66
rect -100 64 -98 69
rect -90 64 -88 69
rect -176 42 -170 44
rect -196 38 -190 40
rect -196 36 -194 38
rect -192 36 -190 38
rect -196 34 -190 36
rect -186 38 -180 40
rect -186 36 -184 38
rect -182 36 -180 38
rect -186 34 -180 36
rect -196 29 -194 34
rect -183 29 -181 34
rect -176 29 -174 42
rect -152 40 -150 44
rect -142 40 -140 51
rect -132 48 -130 51
rect -132 46 -126 48
rect -132 44 -130 46
rect -128 44 -126 46
rect -69 62 -67 66
rect -59 64 -57 69
rect -49 64 -47 69
rect -132 42 -126 44
rect -152 38 -146 40
rect -152 36 -150 38
rect -148 36 -146 38
rect -152 34 -146 36
rect -142 38 -136 40
rect -142 36 -140 38
rect -138 36 -136 38
rect -142 34 -136 36
rect -152 29 -150 34
rect -139 29 -137 34
rect -132 29 -130 42
rect -110 40 -108 44
rect -100 40 -98 51
rect -90 48 -88 51
rect -90 46 -84 48
rect -90 44 -88 46
rect -86 44 -84 46
rect -26 62 -24 66
rect -16 64 -14 69
rect -6 64 -4 69
rect -90 42 -84 44
rect -110 38 -104 40
rect -110 36 -108 38
rect -106 36 -104 38
rect -110 34 -104 36
rect -100 38 -94 40
rect -100 36 -98 38
rect -96 36 -94 38
rect -100 34 -94 36
rect -110 29 -108 34
rect -97 29 -95 34
rect -90 29 -88 42
rect -69 40 -67 44
rect -59 40 -57 51
rect -49 48 -47 51
rect -49 46 -43 48
rect -49 44 -47 46
rect -45 44 -43 46
rect 14 62 16 66
rect 24 64 26 69
rect 34 64 36 69
rect -49 42 -43 44
rect -69 38 -63 40
rect -69 36 -67 38
rect -65 36 -63 38
rect -69 34 -63 36
rect -59 38 -53 40
rect -59 36 -57 38
rect -55 36 -53 38
rect -59 34 -53 36
rect -69 29 -67 34
rect -56 29 -54 34
rect -49 29 -47 42
rect -26 40 -24 44
rect -16 40 -14 51
rect -6 48 -4 51
rect -6 46 0 48
rect -6 44 -4 46
rect -2 44 0 46
rect 57 62 59 66
rect 67 64 69 69
rect 77 64 79 69
rect -6 42 0 44
rect -26 38 -20 40
rect -26 36 -24 38
rect -22 36 -20 38
rect -26 34 -20 36
rect -16 38 -10 40
rect -16 36 -14 38
rect -12 36 -10 38
rect -16 34 -10 36
rect -26 29 -24 34
rect -13 29 -11 34
rect -6 29 -4 42
rect 14 40 16 44
rect 24 40 26 51
rect 34 48 36 51
rect 34 46 40 48
rect 34 44 36 46
rect 38 44 40 46
rect 34 42 40 44
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 29 16 34
rect 27 29 29 34
rect 34 29 36 42
rect 57 40 59 44
rect 67 40 69 51
rect 77 48 79 51
rect 77 46 83 48
rect 77 44 79 46
rect 81 44 83 46
rect 77 42 83 44
rect 57 38 63 40
rect 57 36 59 38
rect 61 36 63 38
rect 57 34 63 36
rect 67 38 73 40
rect 67 36 69 38
rect 71 36 73 38
rect 67 34 73 36
rect 57 29 59 34
rect 70 29 72 34
rect 77 29 79 42
rect -538 16 -536 20
rect -525 13 -523 18
rect -518 13 -516 18
rect -498 16 -496 20
rect -485 13 -483 18
rect -478 13 -476 18
rect -455 16 -453 20
rect -442 13 -440 18
rect -435 13 -433 18
rect -351 16 -349 20
rect -338 13 -336 18
rect -331 13 -329 18
rect -309 16 -307 20
rect -296 13 -294 18
rect -289 13 -287 18
rect -265 16 -263 20
rect -252 13 -250 18
rect -245 13 -243 18
rect -196 16 -194 20
rect -183 13 -181 18
rect -176 13 -174 18
rect -152 16 -150 20
rect -139 13 -137 18
rect -132 13 -130 18
rect -110 16 -108 20
rect -97 13 -95 18
rect -90 13 -88 18
rect -69 16 -67 20
rect -56 13 -54 18
rect -49 13 -47 18
rect -26 16 -24 20
rect -13 13 -11 18
rect -6 13 -4 18
rect 14 16 16 20
rect 27 13 29 18
rect 34 13 36 18
rect 57 16 59 20
rect 70 13 72 18
rect 77 13 79 18
rect -565 0 -563 4
rect -554 0 -552 4
rect -547 0 -545 4
rect -565 -23 -563 -14
rect -527 -6 -525 -1
rect -517 -6 -515 -1
rect -507 -3 -505 2
rect -497 0 -495 4
rect -450 -6 -448 -1
rect -431 1 -409 3
rect -474 -11 -472 -6
rect -554 -23 -552 -20
rect -547 -23 -545 -20
rect -527 -23 -525 -20
rect -517 -23 -515 -20
rect -567 -25 -561 -23
rect -567 -27 -565 -25
rect -563 -27 -561 -25
rect -567 -29 -561 -27
rect -557 -25 -551 -23
rect -557 -27 -555 -25
rect -553 -27 -551 -25
rect -557 -29 -551 -27
rect -547 -25 -525 -23
rect -547 -27 -545 -25
rect -543 -27 -538 -25
rect -536 -27 -525 -25
rect -547 -29 -525 -27
rect -521 -25 -515 -23
rect -521 -27 -519 -25
rect -517 -27 -515 -25
rect -521 -29 -515 -27
rect -507 -26 -505 -13
rect -497 -16 -495 -13
rect -501 -18 -495 -16
rect -501 -20 -499 -18
rect -497 -20 -495 -18
rect -438 -8 -436 -3
rect -431 -8 -429 1
rect -421 -8 -419 -3
rect -411 -8 -409 1
rect -384 -1 -382 4
rect -377 -1 -375 4
rect -367 2 -343 4
rect -367 -1 -365 2
rect -501 -22 -495 -20
rect -507 -28 -501 -26
rect -565 -32 -563 -29
rect -555 -32 -553 -29
rect -545 -32 -543 -29
rect -527 -32 -525 -29
rect -520 -32 -518 -29
rect -507 -30 -505 -28
rect -503 -30 -501 -28
rect -510 -32 -501 -30
rect -510 -35 -508 -32
rect -497 -35 -495 -22
rect -474 -23 -472 -20
rect -450 -23 -448 -18
rect -357 -6 -355 -2
rect -345 -3 -343 2
rect -322 -1 -320 4
rect -315 -1 -313 4
rect -305 2 -282 4
rect -305 -1 -303 2
rect -438 -23 -436 -20
rect -431 -23 -429 -20
rect -421 -23 -419 -20
rect -411 -23 -409 -20
rect -384 -23 -382 -14
rect -377 -17 -375 -14
rect -377 -19 -373 -17
rect -367 -19 -365 -14
rect -295 -6 -293 -2
rect -345 -17 -343 -14
rect -345 -19 -339 -17
rect -375 -23 -373 -19
rect -474 -25 -468 -23
rect -474 -27 -472 -25
rect -470 -27 -468 -25
rect -474 -29 -468 -27
rect -450 -25 -435 -23
rect -450 -27 -448 -25
rect -446 -27 -435 -25
rect -431 -26 -428 -23
rect -450 -29 -435 -27
rect -474 -32 -472 -29
rect -447 -32 -445 -29
rect -437 -32 -435 -29
rect -430 -32 -428 -26
rect -424 -25 -418 -23
rect -424 -27 -422 -25
rect -420 -27 -418 -25
rect -424 -29 -418 -27
rect -411 -25 -404 -23
rect -411 -27 -408 -25
rect -406 -27 -404 -25
rect -411 -29 -404 -27
rect -385 -25 -379 -23
rect -385 -27 -383 -25
rect -381 -27 -379 -25
rect -385 -29 -379 -27
rect -375 -25 -369 -23
rect -375 -27 -373 -25
rect -371 -27 -369 -25
rect -357 -27 -355 -19
rect -345 -21 -343 -19
rect -341 -21 -339 -19
rect -345 -23 -339 -21
rect -322 -23 -320 -14
rect -315 -23 -313 -14
rect -305 -19 -303 -14
rect -284 -9 -282 2
rect -232 -6 -230 -1
rect -213 1 -191 3
rect -295 -22 -293 -19
rect -256 -11 -254 -6
rect -220 -8 -218 -3
rect -213 -8 -211 1
rect -203 -8 -201 -3
rect -193 -8 -191 1
rect -166 -1 -164 4
rect -159 -1 -157 4
rect -149 2 -125 4
rect -149 -1 -147 2
rect -335 -25 -329 -23
rect -335 -27 -333 -25
rect -331 -27 -329 -25
rect -375 -29 -369 -27
rect -365 -29 -329 -27
rect -325 -25 -319 -23
rect -325 -27 -323 -25
rect -321 -27 -319 -25
rect -325 -29 -319 -27
rect -315 -25 -309 -23
rect -315 -27 -313 -25
rect -311 -27 -309 -25
rect -297 -24 -291 -22
rect -297 -26 -295 -24
rect -293 -26 -291 -24
rect -315 -29 -309 -27
rect -305 -28 -291 -26
rect -420 -32 -418 -29
rect -410 -32 -408 -29
rect -385 -32 -383 -29
rect -375 -32 -373 -29
rect -365 -32 -363 -29
rect -325 -32 -323 -29
rect -315 -32 -313 -29
rect -305 -32 -303 -28
rect -510 -53 -508 -48
rect -565 -64 -563 -60
rect -555 -64 -553 -60
rect -545 -64 -543 -60
rect -527 -62 -525 -57
rect -520 -62 -518 -57
rect -474 -55 -472 -50
rect -497 -64 -495 -60
rect -447 -64 -445 -59
rect -437 -64 -435 -59
rect -430 -64 -428 -59
rect -420 -64 -418 -59
rect -410 -64 -408 -59
rect -349 -39 -343 -37
rect -349 -41 -347 -39
rect -345 -41 -343 -39
rect -355 -43 -343 -41
rect -355 -46 -353 -43
rect -345 -46 -343 -43
rect -284 -34 -282 -20
rect -256 -23 -254 -20
rect -232 -23 -230 -18
rect -139 -6 -137 -2
rect -127 -3 -125 2
rect -104 -1 -102 4
rect -97 -1 -95 4
rect -87 2 -64 4
rect -87 -1 -85 2
rect -220 -23 -218 -20
rect -213 -23 -211 -20
rect -203 -23 -201 -20
rect -193 -23 -191 -20
rect -166 -23 -164 -14
rect -159 -17 -157 -14
rect -159 -19 -155 -17
rect -149 -19 -147 -14
rect -77 -6 -75 -2
rect -127 -17 -125 -14
rect -127 -19 -121 -17
rect -157 -23 -155 -19
rect -256 -25 -250 -23
rect -256 -27 -254 -25
rect -252 -27 -250 -25
rect -256 -29 -250 -27
rect -232 -25 -217 -23
rect -232 -27 -230 -25
rect -228 -27 -217 -25
rect -213 -26 -210 -23
rect -232 -29 -217 -27
rect -274 -32 -268 -30
rect -256 -32 -254 -29
rect -229 -32 -227 -29
rect -219 -32 -217 -29
rect -212 -32 -210 -26
rect -206 -25 -200 -23
rect -206 -27 -204 -25
rect -202 -27 -200 -25
rect -206 -29 -200 -27
rect -193 -25 -186 -23
rect -193 -27 -190 -25
rect -188 -27 -186 -25
rect -193 -29 -186 -27
rect -167 -25 -161 -23
rect -167 -27 -165 -25
rect -163 -27 -161 -25
rect -167 -29 -161 -27
rect -157 -25 -151 -23
rect -157 -27 -155 -25
rect -153 -27 -151 -25
rect -139 -27 -137 -19
rect -127 -21 -125 -19
rect -123 -21 -121 -19
rect -127 -23 -121 -21
rect -104 -23 -102 -14
rect -97 -23 -95 -14
rect -87 -19 -85 -14
rect -66 -9 -64 2
rect -27 0 -25 4
rect -16 0 -14 4
rect -9 0 -7 4
rect -77 -22 -75 -19
rect -117 -25 -111 -23
rect -117 -27 -115 -25
rect -113 -27 -111 -25
rect -157 -29 -151 -27
rect -147 -29 -111 -27
rect -107 -25 -101 -23
rect -107 -27 -105 -25
rect -103 -27 -101 -25
rect -107 -29 -101 -27
rect -97 -25 -91 -23
rect -97 -27 -95 -25
rect -93 -27 -91 -25
rect -79 -24 -73 -22
rect -79 -26 -77 -24
rect -75 -26 -73 -24
rect -97 -29 -91 -27
rect -87 -28 -73 -26
rect -202 -32 -200 -29
rect -192 -32 -190 -29
rect -167 -32 -165 -29
rect -157 -32 -155 -29
rect -147 -32 -145 -29
rect -107 -32 -105 -29
rect -97 -32 -95 -29
rect -87 -32 -85 -28
rect -274 -34 -272 -32
rect -270 -34 -268 -32
rect -294 -36 -268 -34
rect -294 -39 -292 -36
rect -284 -39 -282 -36
rect -294 -57 -292 -53
rect -284 -57 -282 -53
rect -256 -55 -254 -50
rect -385 -64 -383 -60
rect -375 -64 -373 -60
rect -365 -64 -363 -60
rect -355 -64 -353 -60
rect -345 -64 -343 -60
rect -325 -64 -323 -60
rect -315 -64 -313 -60
rect -305 -64 -303 -60
rect -229 -64 -227 -59
rect -219 -64 -217 -59
rect -212 -64 -210 -59
rect -202 -64 -200 -59
rect -192 -64 -190 -59
rect -131 -39 -125 -37
rect -131 -41 -129 -39
rect -127 -41 -125 -39
rect -137 -43 -125 -41
rect -137 -46 -135 -43
rect -127 -46 -125 -43
rect -66 -34 -64 -20
rect -27 -23 -25 -14
rect 11 -6 13 -1
rect 21 -6 23 -1
rect 31 -3 33 2
rect 41 0 43 4
rect -16 -23 -14 -20
rect -9 -23 -7 -20
rect 11 -23 13 -20
rect 21 -23 23 -20
rect -29 -25 -23 -23
rect -29 -27 -27 -25
rect -25 -27 -23 -25
rect -29 -29 -23 -27
rect -19 -25 -13 -23
rect -19 -27 -17 -25
rect -15 -27 -13 -25
rect -19 -29 -13 -27
rect -9 -25 13 -23
rect -9 -27 -7 -25
rect -5 -27 0 -25
rect 2 -27 13 -25
rect -9 -29 13 -27
rect 17 -25 23 -23
rect 17 -27 19 -25
rect 21 -27 23 -25
rect 17 -29 23 -27
rect 31 -26 33 -13
rect 41 -16 43 -13
rect 37 -18 43 -16
rect 37 -20 39 -18
rect 41 -20 43 -18
rect 37 -22 43 -20
rect 31 -28 37 -26
rect -56 -32 -50 -30
rect -27 -32 -25 -29
rect -17 -32 -15 -29
rect -7 -32 -5 -29
rect 11 -32 13 -29
rect 18 -32 20 -29
rect 31 -30 33 -28
rect 35 -30 37 -28
rect 28 -32 37 -30
rect -56 -34 -54 -32
rect -52 -34 -50 -32
rect -76 -36 -50 -34
rect -76 -39 -74 -36
rect -66 -39 -64 -36
rect -76 -57 -74 -53
rect -66 -57 -64 -53
rect -167 -64 -165 -60
rect -157 -64 -155 -60
rect -147 -64 -145 -60
rect -137 -64 -135 -60
rect -127 -64 -125 -60
rect -107 -64 -105 -60
rect -97 -64 -95 -60
rect -87 -64 -85 -60
rect 28 -35 30 -32
rect 41 -35 43 -22
rect 28 -53 30 -48
rect -27 -64 -25 -60
rect -17 -64 -15 -60
rect -7 -64 -5 -60
rect 11 -62 13 -57
rect 18 -62 20 -57
rect 41 -64 43 -60
rect -483 -73 -481 -68
rect -473 -73 -471 -68
rect -466 -73 -464 -68
rect -456 -73 -454 -68
rect -446 -73 -444 -68
rect -421 -72 -419 -68
rect -411 -72 -409 -68
rect -401 -72 -399 -68
rect -391 -72 -389 -68
rect -381 -72 -379 -68
rect -361 -72 -359 -68
rect -351 -72 -349 -68
rect -341 -72 -339 -68
rect -510 -82 -508 -77
rect -391 -89 -389 -86
rect -381 -89 -379 -86
rect -391 -91 -379 -89
rect -385 -93 -383 -91
rect -381 -93 -379 -91
rect -385 -95 -379 -93
rect -263 -73 -261 -68
rect -253 -73 -251 -68
rect -246 -73 -244 -68
rect -236 -73 -234 -68
rect -226 -73 -224 -68
rect -201 -72 -199 -68
rect -191 -72 -189 -68
rect -181 -72 -179 -68
rect -171 -72 -169 -68
rect -161 -72 -159 -68
rect -141 -72 -139 -68
rect -131 -72 -129 -68
rect -121 -72 -119 -68
rect -330 -79 -328 -75
rect -320 -79 -318 -75
rect -290 -82 -288 -77
rect -330 -96 -328 -93
rect -320 -96 -318 -93
rect -330 -98 -304 -96
rect -510 -103 -508 -100
rect -483 -103 -481 -100
rect -473 -103 -471 -100
rect -510 -105 -504 -103
rect -510 -107 -508 -105
rect -506 -107 -504 -105
rect -510 -109 -504 -107
rect -486 -105 -471 -103
rect -486 -107 -484 -105
rect -482 -107 -471 -105
rect -466 -106 -464 -100
rect -456 -103 -454 -100
rect -446 -103 -444 -100
rect -421 -103 -419 -100
rect -411 -103 -409 -100
rect -401 -103 -399 -100
rect -361 -103 -359 -100
rect -351 -103 -349 -100
rect -486 -109 -471 -107
rect -467 -109 -464 -106
rect -460 -105 -454 -103
rect -460 -107 -458 -105
rect -456 -107 -454 -105
rect -460 -109 -454 -107
rect -447 -105 -440 -103
rect -447 -107 -444 -105
rect -442 -107 -440 -105
rect -447 -109 -440 -107
rect -421 -105 -415 -103
rect -421 -107 -419 -105
rect -417 -107 -415 -105
rect -421 -109 -415 -107
rect -411 -105 -405 -103
rect -401 -105 -365 -103
rect -411 -107 -409 -105
rect -407 -107 -405 -105
rect -411 -109 -405 -107
rect -510 -112 -508 -109
rect -486 -114 -484 -109
rect -474 -112 -472 -109
rect -467 -112 -465 -109
rect -457 -112 -455 -109
rect -447 -112 -445 -109
rect -510 -126 -508 -121
rect -420 -118 -418 -109
rect -411 -113 -409 -109
rect -393 -113 -391 -105
rect -371 -107 -369 -105
rect -367 -107 -365 -105
rect -371 -109 -365 -107
rect -361 -105 -355 -103
rect -361 -107 -359 -105
rect -357 -107 -355 -105
rect -361 -109 -355 -107
rect -351 -105 -345 -103
rect -351 -107 -349 -105
rect -347 -107 -345 -105
rect -341 -104 -339 -100
rect -341 -106 -327 -104
rect -351 -109 -345 -107
rect -333 -108 -331 -106
rect -329 -108 -327 -106
rect -381 -111 -375 -109
rect -381 -113 -379 -111
rect -377 -113 -375 -111
rect -413 -115 -409 -113
rect -413 -118 -411 -115
rect -403 -118 -401 -113
rect -486 -131 -484 -126
rect -474 -129 -472 -124
rect -467 -133 -465 -124
rect -457 -129 -455 -124
rect -447 -133 -445 -124
rect -467 -135 -445 -133
rect -381 -115 -375 -113
rect -381 -118 -379 -115
rect -358 -118 -356 -109
rect -351 -118 -349 -109
rect -333 -110 -327 -108
rect -331 -113 -329 -110
rect -320 -112 -318 -98
rect -310 -100 -308 -98
rect -306 -100 -304 -98
rect -171 -89 -169 -86
rect -161 -89 -159 -86
rect -171 -91 -159 -89
rect -165 -93 -163 -91
rect -161 -93 -159 -91
rect -165 -95 -159 -93
rect -68 -72 -66 -68
rect -58 -72 -56 -68
rect -48 -72 -46 -68
rect -110 -79 -108 -75
rect -100 -79 -98 -75
rect -110 -96 -108 -93
rect -100 -96 -98 -93
rect -110 -98 -84 -96
rect -310 -102 -304 -100
rect -290 -103 -288 -100
rect -263 -103 -261 -100
rect -253 -103 -251 -100
rect -290 -105 -284 -103
rect -290 -107 -288 -105
rect -286 -107 -284 -105
rect -290 -109 -284 -107
rect -266 -105 -251 -103
rect -266 -107 -264 -105
rect -262 -107 -251 -105
rect -246 -106 -244 -100
rect -236 -103 -234 -100
rect -226 -103 -224 -100
rect -201 -103 -199 -100
rect -191 -103 -189 -100
rect -181 -103 -179 -100
rect -141 -103 -139 -100
rect -131 -103 -129 -100
rect -266 -109 -251 -107
rect -247 -109 -244 -106
rect -240 -105 -234 -103
rect -240 -107 -238 -105
rect -236 -107 -234 -105
rect -240 -109 -234 -107
rect -227 -105 -220 -103
rect -227 -107 -224 -105
rect -222 -107 -220 -105
rect -227 -109 -220 -107
rect -201 -105 -195 -103
rect -201 -107 -199 -105
rect -197 -107 -195 -105
rect -201 -109 -195 -107
rect -191 -105 -185 -103
rect -181 -105 -145 -103
rect -191 -107 -189 -105
rect -187 -107 -185 -105
rect -191 -109 -185 -107
rect -290 -112 -288 -109
rect -341 -118 -339 -113
rect -393 -130 -391 -126
rect -420 -136 -418 -131
rect -413 -136 -411 -131
rect -403 -134 -401 -131
rect -381 -134 -379 -129
rect -403 -136 -379 -134
rect -266 -114 -264 -109
rect -254 -112 -252 -109
rect -247 -112 -245 -109
rect -237 -112 -235 -109
rect -227 -112 -225 -109
rect -331 -130 -329 -126
rect -358 -136 -356 -131
rect -351 -136 -349 -131
rect -341 -134 -339 -131
rect -320 -134 -318 -123
rect -290 -126 -288 -121
rect -200 -118 -198 -109
rect -191 -113 -189 -109
rect -173 -113 -171 -105
rect -151 -107 -149 -105
rect -147 -107 -145 -105
rect -151 -109 -145 -107
rect -141 -105 -135 -103
rect -141 -107 -139 -105
rect -137 -107 -135 -105
rect -141 -109 -135 -107
rect -131 -105 -125 -103
rect -131 -107 -129 -105
rect -127 -107 -125 -105
rect -121 -104 -119 -100
rect -121 -106 -107 -104
rect -131 -109 -125 -107
rect -113 -108 -111 -106
rect -109 -108 -107 -106
rect -161 -111 -155 -109
rect -161 -113 -159 -111
rect -157 -113 -155 -111
rect -193 -115 -189 -113
rect -193 -118 -191 -115
rect -183 -118 -181 -113
rect -341 -136 -318 -134
rect -266 -131 -264 -126
rect -254 -129 -252 -124
rect -247 -133 -245 -124
rect -237 -129 -235 -124
rect -227 -133 -225 -124
rect -247 -135 -225 -133
rect -161 -115 -155 -113
rect -161 -118 -159 -115
rect -138 -118 -136 -109
rect -131 -118 -129 -109
rect -113 -110 -107 -108
rect -111 -113 -109 -110
rect -100 -112 -98 -98
rect -90 -100 -88 -98
rect -86 -100 -84 -98
rect -30 -75 -28 -70
rect -23 -75 -21 -70
rect 0 -72 2 -68
rect -13 -84 -11 -79
rect -13 -100 -11 -97
rect -90 -102 -84 -100
rect -68 -103 -66 -100
rect -58 -103 -56 -100
rect -48 -103 -46 -100
rect -30 -103 -28 -100
rect -23 -103 -21 -100
rect -13 -102 -4 -100
rect -70 -105 -64 -103
rect -70 -107 -68 -105
rect -66 -107 -64 -105
rect -70 -109 -64 -107
rect -60 -105 -54 -103
rect -60 -107 -58 -105
rect -56 -107 -54 -105
rect -60 -109 -54 -107
rect -50 -105 -28 -103
rect -50 -107 -48 -105
rect -46 -107 -41 -105
rect -39 -107 -28 -105
rect -50 -109 -28 -107
rect -24 -105 -18 -103
rect -24 -107 -22 -105
rect -20 -107 -18 -105
rect -24 -109 -18 -107
rect -121 -118 -119 -113
rect -173 -130 -171 -126
rect -200 -136 -198 -131
rect -193 -136 -191 -131
rect -183 -134 -181 -131
rect -161 -134 -159 -129
rect -183 -136 -159 -134
rect -68 -118 -66 -109
rect -57 -112 -55 -109
rect -50 -112 -48 -109
rect -30 -112 -28 -109
rect -20 -112 -18 -109
rect -10 -104 -8 -102
rect -6 -104 -4 -102
rect -10 -106 -4 -104
rect -111 -130 -109 -126
rect -138 -136 -136 -131
rect -131 -136 -129 -131
rect -121 -134 -119 -131
rect -100 -134 -98 -123
rect -121 -136 -98 -134
rect -10 -119 -8 -106
rect 0 -110 2 -97
rect -4 -112 2 -110
rect -4 -114 -2 -112
rect 0 -114 2 -112
rect -4 -116 2 -114
rect 0 -119 2 -116
rect -30 -131 -28 -126
rect -20 -131 -18 -126
rect -68 -136 -66 -132
rect -57 -136 -55 -132
rect -50 -136 -48 -132
rect -10 -134 -8 -129
rect 0 -136 2 -132
<< ndif >>
rect -543 26 -538 29
rect -545 24 -538 26
rect -545 22 -543 24
rect -541 22 -538 24
rect -545 20 -538 22
rect -536 20 -525 29
rect -534 18 -525 20
rect -523 18 -518 29
rect -516 24 -511 29
rect -503 26 -498 29
rect -505 24 -498 26
rect -516 22 -509 24
rect -516 20 -513 22
rect -511 20 -509 22
rect -505 22 -503 24
rect -501 22 -498 24
rect -505 20 -498 22
rect -496 20 -485 29
rect -516 18 -509 20
rect -534 12 -527 18
rect -494 18 -485 20
rect -483 18 -478 29
rect -476 24 -471 29
rect -460 26 -455 29
rect -462 24 -455 26
rect -476 22 -469 24
rect -476 20 -473 22
rect -471 20 -469 22
rect -462 22 -460 24
rect -458 22 -455 24
rect -462 20 -455 22
rect -453 20 -442 29
rect -476 18 -469 20
rect -534 10 -532 12
rect -530 10 -527 12
rect -534 8 -527 10
rect -494 12 -487 18
rect -451 18 -442 20
rect -440 18 -435 29
rect -433 24 -428 29
rect -356 26 -351 29
rect -358 24 -351 26
rect -433 22 -426 24
rect -433 20 -430 22
rect -428 20 -426 22
rect -358 22 -356 24
rect -354 22 -351 24
rect -358 20 -351 22
rect -349 20 -338 29
rect -433 18 -426 20
rect -494 10 -492 12
rect -490 10 -487 12
rect -494 8 -487 10
rect -451 12 -444 18
rect -347 18 -338 20
rect -336 18 -331 29
rect -329 24 -324 29
rect -314 26 -309 29
rect -316 24 -309 26
rect -329 22 -322 24
rect -329 20 -326 22
rect -324 20 -322 22
rect -316 22 -314 24
rect -312 22 -309 24
rect -316 20 -309 22
rect -307 20 -296 29
rect -329 18 -322 20
rect -451 10 -449 12
rect -447 10 -444 12
rect -451 8 -444 10
rect -347 12 -340 18
rect -305 18 -296 20
rect -294 18 -289 29
rect -287 24 -282 29
rect -270 26 -265 29
rect -272 24 -265 26
rect -287 22 -280 24
rect -287 20 -284 22
rect -282 20 -280 22
rect -272 22 -270 24
rect -268 22 -265 24
rect -272 20 -265 22
rect -263 20 -252 29
rect -287 18 -280 20
rect -347 10 -345 12
rect -343 10 -340 12
rect -347 8 -340 10
rect -305 12 -298 18
rect -261 18 -252 20
rect -250 18 -245 29
rect -243 24 -238 29
rect -201 26 -196 29
rect -203 24 -196 26
rect -243 22 -236 24
rect -243 20 -240 22
rect -238 20 -236 22
rect -203 22 -201 24
rect -199 22 -196 24
rect -203 20 -196 22
rect -194 20 -183 29
rect -243 18 -236 20
rect -305 10 -303 12
rect -301 10 -298 12
rect -305 8 -298 10
rect -261 12 -254 18
rect -192 18 -183 20
rect -181 18 -176 29
rect -174 24 -169 29
rect -157 26 -152 29
rect -159 24 -152 26
rect -174 22 -167 24
rect -174 20 -171 22
rect -169 20 -167 22
rect -159 22 -157 24
rect -155 22 -152 24
rect -159 20 -152 22
rect -150 20 -139 29
rect -174 18 -167 20
rect -261 10 -259 12
rect -257 10 -254 12
rect -261 8 -254 10
rect -192 12 -185 18
rect -148 18 -139 20
rect -137 18 -132 29
rect -130 24 -125 29
rect -115 26 -110 29
rect -117 24 -110 26
rect -130 22 -123 24
rect -130 20 -127 22
rect -125 20 -123 22
rect -117 22 -115 24
rect -113 22 -110 24
rect -117 20 -110 22
rect -108 20 -97 29
rect -130 18 -123 20
rect -192 10 -190 12
rect -188 10 -185 12
rect -192 8 -185 10
rect -148 12 -141 18
rect -106 18 -97 20
rect -95 18 -90 29
rect -88 24 -83 29
rect -74 26 -69 29
rect -76 24 -69 26
rect -88 22 -81 24
rect -88 20 -85 22
rect -83 20 -81 22
rect -76 22 -74 24
rect -72 22 -69 24
rect -76 20 -69 22
rect -67 20 -56 29
rect -88 18 -81 20
rect -148 10 -146 12
rect -144 10 -141 12
rect -148 8 -141 10
rect -106 12 -99 18
rect -65 18 -56 20
rect -54 18 -49 29
rect -47 24 -42 29
rect -31 26 -26 29
rect -33 24 -26 26
rect -47 22 -40 24
rect -47 20 -44 22
rect -42 20 -40 22
rect -33 22 -31 24
rect -29 22 -26 24
rect -33 20 -26 22
rect -24 20 -13 29
rect -47 18 -40 20
rect -106 10 -104 12
rect -102 10 -99 12
rect -106 8 -99 10
rect -65 12 -58 18
rect -22 18 -13 20
rect -11 18 -6 29
rect -4 24 1 29
rect 9 26 14 29
rect 7 24 14 26
rect -4 22 3 24
rect -4 20 -1 22
rect 1 20 3 22
rect 7 22 9 24
rect 11 22 14 24
rect 7 20 14 22
rect 16 20 27 29
rect -4 18 3 20
rect -65 10 -63 12
rect -61 10 -58 12
rect -65 8 -58 10
rect -22 12 -15 18
rect 18 18 27 20
rect 29 18 34 29
rect 36 24 41 29
rect 52 26 57 29
rect 50 24 57 26
rect 36 22 43 24
rect 36 20 39 22
rect 41 20 43 22
rect 50 22 52 24
rect 54 22 57 24
rect 50 20 57 22
rect 59 20 70 29
rect 36 18 43 20
rect -22 10 -20 12
rect -18 10 -15 12
rect -22 8 -15 10
rect 18 12 25 18
rect 61 18 70 20
rect 72 18 77 29
rect 79 24 84 29
rect 79 22 86 24
rect 79 20 82 22
rect 84 20 86 22
rect 79 18 86 20
rect 18 10 20 12
rect 22 10 25 12
rect 18 8 25 10
rect 61 12 68 18
rect 61 10 63 12
rect 65 10 68 12
rect 61 8 68 10
rect -570 -7 -565 0
rect -572 -9 -565 -7
rect -572 -11 -570 -9
rect -568 -11 -565 -9
rect -572 -14 -565 -11
rect -563 -2 -554 0
rect -563 -4 -559 -2
rect -557 -4 -554 -2
rect -563 -14 -554 -4
rect -561 -20 -554 -14
rect -552 -20 -547 0
rect -545 -7 -540 0
rect -502 -3 -497 0
rect -512 -6 -507 -3
rect -545 -9 -538 -7
rect -545 -11 -542 -9
rect -540 -11 -538 -9
rect -545 -13 -538 -11
rect -534 -9 -527 -6
rect -534 -11 -532 -9
rect -530 -11 -527 -9
rect -545 -20 -540 -13
rect -534 -16 -527 -11
rect -534 -18 -532 -16
rect -530 -18 -527 -16
rect -534 -20 -527 -18
rect -525 -16 -517 -6
rect -525 -18 -522 -16
rect -520 -18 -517 -16
rect -525 -20 -517 -18
rect -515 -8 -507 -6
rect -515 -10 -512 -8
rect -510 -10 -507 -8
rect -515 -13 -507 -10
rect -505 -5 -497 -3
rect -505 -7 -502 -5
rect -500 -7 -497 -5
rect -505 -13 -497 -7
rect -495 -7 -490 0
rect -446 1 -440 3
rect -446 -1 -444 1
rect -442 -1 -440 1
rect -446 -6 -440 -1
rect -495 -9 -488 -7
rect -495 -11 -492 -9
rect -490 -11 -488 -9
rect -457 -8 -450 -6
rect -457 -10 -455 -8
rect -453 -10 -450 -8
rect -495 -13 -488 -11
rect -515 -20 -510 -13
rect -479 -14 -474 -11
rect -481 -16 -474 -14
rect -481 -18 -479 -16
rect -477 -18 -474 -16
rect -481 -20 -474 -18
rect -472 -13 -461 -11
rect -457 -12 -450 -10
rect -472 -15 -465 -13
rect -463 -15 -461 -13
rect -472 -20 -461 -15
rect -455 -18 -450 -12
rect -448 -8 -440 -6
rect -392 1 -386 3
rect -392 -1 -390 1
rect -388 -1 -386 1
rect -448 -18 -438 -8
rect -446 -20 -438 -18
rect -436 -20 -431 -8
rect -429 -16 -421 -8
rect -429 -18 -426 -16
rect -424 -18 -421 -16
rect -429 -20 -421 -18
rect -419 -10 -411 -8
rect -419 -12 -416 -10
rect -414 -12 -411 -10
rect -419 -20 -411 -12
rect -409 -10 -401 -8
rect -409 -12 -406 -10
rect -404 -12 -401 -10
rect -409 -20 -401 -12
rect -392 -14 -384 -1
rect -382 -14 -377 -1
rect -375 -9 -367 -1
rect -375 -11 -372 -9
rect -370 -11 -367 -9
rect -375 -14 -367 -11
rect -365 -6 -360 -1
rect -353 -2 -347 0
rect -353 -4 -351 -2
rect -349 -3 -347 -2
rect -330 1 -324 3
rect -330 -1 -328 1
rect -326 -1 -324 1
rect -349 -4 -345 -3
rect -353 -6 -345 -4
rect -365 -10 -357 -6
rect -365 -12 -362 -10
rect -360 -12 -357 -10
rect -365 -14 -357 -12
rect -362 -19 -357 -14
rect -355 -14 -345 -6
rect -343 -8 -338 -3
rect -343 -10 -336 -8
rect -343 -12 -340 -10
rect -338 -12 -336 -10
rect -343 -14 -336 -12
rect -330 -14 -322 -1
rect -320 -14 -315 -1
rect -313 -9 -305 -1
rect -313 -11 -310 -9
rect -308 -11 -305 -9
rect -313 -14 -305 -11
rect -303 -6 -298 -1
rect -303 -10 -295 -6
rect -303 -12 -300 -10
rect -298 -12 -295 -10
rect -303 -14 -295 -12
rect -355 -19 -347 -14
rect -300 -19 -295 -14
rect -293 -8 -286 -6
rect -293 -10 -290 -8
rect -288 -9 -286 -8
rect -228 1 -222 3
rect -228 -1 -226 1
rect -224 -1 -222 1
rect -228 -6 -222 -1
rect -288 -10 -284 -9
rect -293 -19 -284 -10
rect -289 -20 -284 -19
rect -282 -14 -277 -9
rect -239 -8 -232 -6
rect -239 -10 -237 -8
rect -235 -10 -232 -8
rect -261 -14 -256 -11
rect -282 -16 -275 -14
rect -282 -18 -279 -16
rect -277 -18 -275 -16
rect -282 -20 -275 -18
rect -263 -16 -256 -14
rect -263 -18 -261 -16
rect -259 -18 -256 -16
rect -263 -20 -256 -18
rect -254 -13 -243 -11
rect -239 -12 -232 -10
rect -254 -15 -247 -13
rect -245 -15 -243 -13
rect -254 -20 -243 -15
rect -237 -18 -232 -12
rect -230 -8 -222 -6
rect -174 1 -168 3
rect -174 -1 -172 1
rect -170 -1 -168 1
rect -230 -18 -220 -8
rect -228 -20 -220 -18
rect -218 -20 -213 -8
rect -211 -16 -203 -8
rect -211 -18 -208 -16
rect -206 -18 -203 -16
rect -211 -20 -203 -18
rect -201 -10 -193 -8
rect -201 -12 -198 -10
rect -196 -12 -193 -10
rect -201 -20 -193 -12
rect -191 -10 -183 -8
rect -191 -12 -188 -10
rect -186 -12 -183 -10
rect -191 -20 -183 -12
rect -174 -14 -166 -1
rect -164 -14 -159 -1
rect -157 -9 -149 -1
rect -157 -11 -154 -9
rect -152 -11 -149 -9
rect -157 -14 -149 -11
rect -147 -6 -142 -1
rect -135 -2 -129 0
rect -135 -4 -133 -2
rect -131 -3 -129 -2
rect -112 1 -106 3
rect -112 -1 -110 1
rect -108 -1 -106 1
rect -131 -4 -127 -3
rect -135 -6 -127 -4
rect -147 -10 -139 -6
rect -147 -12 -144 -10
rect -142 -12 -139 -10
rect -147 -14 -139 -12
rect -144 -19 -139 -14
rect -137 -14 -127 -6
rect -125 -8 -120 -3
rect -125 -10 -118 -8
rect -125 -12 -122 -10
rect -120 -12 -118 -10
rect -125 -14 -118 -12
rect -112 -14 -104 -1
rect -102 -14 -97 -1
rect -95 -9 -87 -1
rect -95 -11 -92 -9
rect -90 -11 -87 -9
rect -95 -14 -87 -11
rect -85 -6 -80 -1
rect -85 -10 -77 -6
rect -85 -12 -82 -10
rect -80 -12 -77 -10
rect -85 -14 -77 -12
rect -137 -19 -129 -14
rect -82 -19 -77 -14
rect -75 -8 -68 -6
rect -75 -10 -72 -8
rect -70 -9 -68 -8
rect -32 -7 -27 0
rect -34 -9 -27 -7
rect -70 -10 -66 -9
rect -75 -19 -66 -10
rect -71 -20 -66 -19
rect -64 -14 -59 -9
rect -34 -11 -32 -9
rect -30 -11 -27 -9
rect -34 -14 -27 -11
rect -25 -2 -16 0
rect -25 -4 -21 -2
rect -19 -4 -16 -2
rect -25 -14 -16 -4
rect -64 -16 -57 -14
rect -64 -18 -61 -16
rect -59 -18 -57 -16
rect -64 -20 -57 -18
rect -23 -20 -16 -14
rect -14 -20 -9 0
rect -7 -7 -2 0
rect 36 -3 41 0
rect 26 -6 31 -3
rect -7 -9 0 -7
rect -7 -11 -4 -9
rect -2 -11 0 -9
rect -7 -13 0 -11
rect 4 -9 11 -6
rect 4 -11 6 -9
rect 8 -11 11 -9
rect -7 -20 -2 -13
rect 4 -16 11 -11
rect 4 -18 6 -16
rect 8 -18 11 -16
rect 4 -20 11 -18
rect 13 -16 21 -6
rect 13 -18 16 -16
rect 18 -18 21 -16
rect 13 -20 21 -18
rect 23 -8 31 -6
rect 23 -10 26 -8
rect 28 -10 31 -8
rect 23 -13 31 -10
rect 33 -5 41 -3
rect 33 -7 36 -5
rect 38 -7 41 -5
rect 33 -13 41 -7
rect 43 -7 48 0
rect 43 -9 50 -7
rect 43 -11 46 -9
rect 48 -11 50 -9
rect 43 -13 50 -11
rect 23 -20 28 -13
rect -517 -114 -510 -112
rect -517 -116 -515 -114
rect -513 -116 -510 -114
rect -517 -118 -510 -116
rect -515 -121 -510 -118
rect -508 -117 -497 -112
rect -482 -114 -474 -112
rect -508 -119 -501 -117
rect -499 -119 -497 -117
rect -508 -121 -497 -119
rect -491 -120 -486 -114
rect -493 -122 -486 -120
rect -493 -124 -491 -122
rect -489 -124 -486 -122
rect -493 -126 -486 -124
rect -484 -124 -474 -114
rect -472 -124 -467 -112
rect -465 -114 -457 -112
rect -465 -116 -462 -114
rect -460 -116 -457 -114
rect -465 -124 -457 -116
rect -455 -120 -447 -112
rect -455 -122 -452 -120
rect -450 -122 -447 -120
rect -455 -124 -447 -122
rect -445 -120 -437 -112
rect -398 -118 -393 -113
rect -445 -122 -442 -120
rect -440 -122 -437 -120
rect -445 -124 -437 -122
rect -484 -126 -476 -124
rect -482 -131 -476 -126
rect -482 -133 -480 -131
rect -478 -133 -476 -131
rect -482 -135 -476 -133
rect -428 -131 -420 -118
rect -418 -131 -413 -118
rect -411 -121 -403 -118
rect -411 -123 -408 -121
rect -406 -123 -403 -121
rect -411 -131 -403 -123
rect -401 -120 -393 -118
rect -401 -122 -398 -120
rect -396 -122 -393 -120
rect -401 -126 -393 -122
rect -391 -118 -383 -113
rect -325 -113 -320 -112
rect -336 -118 -331 -113
rect -391 -126 -381 -118
rect -401 -131 -396 -126
rect -389 -128 -381 -126
rect -389 -130 -387 -128
rect -385 -129 -381 -128
rect -379 -120 -372 -118
rect -379 -122 -376 -120
rect -374 -122 -372 -120
rect -379 -124 -372 -122
rect -379 -129 -374 -124
rect -385 -130 -383 -129
rect -428 -133 -426 -131
rect -424 -133 -422 -131
rect -428 -135 -422 -133
rect -389 -132 -383 -130
rect -366 -131 -358 -118
rect -356 -131 -351 -118
rect -349 -121 -341 -118
rect -349 -123 -346 -121
rect -344 -123 -341 -121
rect -349 -131 -341 -123
rect -339 -120 -331 -118
rect -339 -122 -336 -120
rect -334 -122 -331 -120
rect -339 -126 -331 -122
rect -329 -122 -320 -113
rect -329 -124 -326 -122
rect -324 -123 -320 -122
rect -318 -114 -311 -112
rect -318 -116 -315 -114
rect -313 -116 -311 -114
rect -318 -118 -311 -116
rect -297 -114 -290 -112
rect -297 -116 -295 -114
rect -293 -116 -290 -114
rect -297 -118 -290 -116
rect -318 -123 -313 -118
rect -295 -121 -290 -118
rect -288 -117 -277 -112
rect -262 -114 -254 -112
rect -288 -119 -281 -117
rect -279 -119 -277 -117
rect -288 -121 -277 -119
rect -271 -120 -266 -114
rect -324 -124 -322 -123
rect -329 -126 -322 -124
rect -339 -131 -334 -126
rect -366 -133 -364 -131
rect -362 -133 -360 -131
rect -366 -135 -360 -133
rect -273 -122 -266 -120
rect -273 -124 -271 -122
rect -269 -124 -266 -122
rect -273 -126 -266 -124
rect -264 -124 -254 -114
rect -252 -124 -247 -112
rect -245 -114 -237 -112
rect -245 -116 -242 -114
rect -240 -116 -237 -114
rect -245 -124 -237 -116
rect -235 -120 -227 -112
rect -235 -122 -232 -120
rect -230 -122 -227 -120
rect -235 -124 -227 -122
rect -225 -120 -217 -112
rect -178 -118 -173 -113
rect -225 -122 -222 -120
rect -220 -122 -217 -120
rect -225 -124 -217 -122
rect -264 -126 -256 -124
rect -262 -131 -256 -126
rect -262 -133 -260 -131
rect -258 -133 -256 -131
rect -262 -135 -256 -133
rect -208 -131 -200 -118
rect -198 -131 -193 -118
rect -191 -121 -183 -118
rect -191 -123 -188 -121
rect -186 -123 -183 -121
rect -191 -131 -183 -123
rect -181 -120 -173 -118
rect -181 -122 -178 -120
rect -176 -122 -173 -120
rect -181 -126 -173 -122
rect -171 -118 -163 -113
rect -105 -113 -100 -112
rect -116 -118 -111 -113
rect -171 -126 -161 -118
rect -181 -131 -176 -126
rect -169 -128 -161 -126
rect -169 -130 -167 -128
rect -165 -129 -161 -128
rect -159 -120 -152 -118
rect -159 -122 -156 -120
rect -154 -122 -152 -120
rect -159 -124 -152 -122
rect -159 -129 -154 -124
rect -165 -130 -163 -129
rect -208 -133 -206 -131
rect -204 -133 -202 -131
rect -208 -135 -202 -133
rect -169 -132 -163 -130
rect -146 -131 -138 -118
rect -136 -131 -131 -118
rect -129 -121 -121 -118
rect -129 -123 -126 -121
rect -124 -123 -121 -121
rect -129 -131 -121 -123
rect -119 -120 -111 -118
rect -119 -122 -116 -120
rect -114 -122 -111 -120
rect -119 -126 -111 -122
rect -109 -122 -100 -113
rect -109 -124 -106 -122
rect -104 -123 -100 -122
rect -98 -114 -91 -112
rect -98 -116 -95 -114
rect -93 -116 -91 -114
rect -98 -118 -91 -116
rect -64 -118 -57 -112
rect -98 -123 -93 -118
rect -75 -121 -68 -118
rect -75 -123 -73 -121
rect -71 -123 -68 -121
rect -104 -124 -102 -123
rect -109 -126 -102 -124
rect -119 -131 -114 -126
rect -146 -133 -144 -131
rect -142 -133 -140 -131
rect -146 -135 -140 -133
rect -75 -125 -68 -123
rect -73 -132 -68 -125
rect -66 -128 -57 -118
rect -66 -130 -62 -128
rect -60 -130 -57 -128
rect -66 -132 -57 -130
rect -55 -132 -50 -112
rect -48 -119 -43 -112
rect -37 -114 -30 -112
rect -37 -116 -35 -114
rect -33 -116 -30 -114
rect -48 -121 -41 -119
rect -48 -123 -45 -121
rect -43 -123 -41 -121
rect -48 -125 -41 -123
rect -37 -121 -30 -116
rect -37 -123 -35 -121
rect -33 -123 -30 -121
rect -48 -132 -43 -125
rect -37 -126 -30 -123
rect -28 -114 -20 -112
rect -28 -116 -25 -114
rect -23 -116 -20 -114
rect -28 -126 -20 -116
rect -18 -119 -13 -112
rect -18 -122 -10 -119
rect -18 -124 -15 -122
rect -13 -124 -10 -122
rect -18 -126 -10 -124
rect -15 -129 -10 -126
rect -8 -125 0 -119
rect -8 -127 -5 -125
rect -3 -127 0 -125
rect -8 -129 0 -127
rect -5 -132 0 -129
rect 2 -121 9 -119
rect 2 -123 5 -121
rect 7 -123 9 -121
rect 2 -125 9 -123
rect 2 -132 7 -125
<< pdif >>
rect -534 62 -528 64
rect -543 57 -538 62
rect -545 55 -538 57
rect -545 53 -543 55
rect -541 53 -538 55
rect -545 48 -538 53
rect -545 46 -543 48
rect -541 46 -538 48
rect -545 44 -538 46
rect -536 60 -528 62
rect -536 58 -533 60
rect -531 58 -528 60
rect -536 51 -528 58
rect -526 62 -518 64
rect -526 60 -523 62
rect -521 60 -518 62
rect -526 55 -518 60
rect -526 53 -523 55
rect -521 53 -518 55
rect -526 51 -518 53
rect -516 62 -509 64
rect -494 62 -488 64
rect -516 60 -513 62
rect -511 60 -509 62
rect -516 51 -509 60
rect -503 57 -498 62
rect -505 55 -498 57
rect -505 53 -503 55
rect -501 53 -498 55
rect -536 44 -530 51
rect -505 48 -498 53
rect -505 46 -503 48
rect -501 46 -498 48
rect -505 44 -498 46
rect -496 60 -488 62
rect -496 58 -493 60
rect -491 58 -488 60
rect -496 51 -488 58
rect -486 62 -478 64
rect -486 60 -483 62
rect -481 60 -478 62
rect -486 55 -478 60
rect -486 53 -483 55
rect -481 53 -478 55
rect -486 51 -478 53
rect -476 62 -469 64
rect -451 62 -445 64
rect -476 60 -473 62
rect -471 60 -469 62
rect -476 51 -469 60
rect -460 57 -455 62
rect -462 55 -455 57
rect -462 53 -460 55
rect -458 53 -455 55
rect -496 44 -490 51
rect -462 48 -455 53
rect -462 46 -460 48
rect -458 46 -455 48
rect -462 44 -455 46
rect -453 60 -445 62
rect -453 58 -450 60
rect -448 58 -445 60
rect -453 51 -445 58
rect -443 62 -435 64
rect -443 60 -440 62
rect -438 60 -435 62
rect -443 55 -435 60
rect -443 53 -440 55
rect -438 53 -435 55
rect -443 51 -435 53
rect -433 62 -426 64
rect -347 62 -341 64
rect -433 60 -430 62
rect -428 60 -426 62
rect -433 51 -426 60
rect -356 57 -351 62
rect -358 55 -351 57
rect -358 53 -356 55
rect -354 53 -351 55
rect -453 44 -447 51
rect -358 48 -351 53
rect -358 46 -356 48
rect -354 46 -351 48
rect -358 44 -351 46
rect -349 60 -341 62
rect -349 58 -346 60
rect -344 58 -341 60
rect -349 51 -341 58
rect -339 62 -331 64
rect -339 60 -336 62
rect -334 60 -331 62
rect -339 55 -331 60
rect -339 53 -336 55
rect -334 53 -331 55
rect -339 51 -331 53
rect -329 62 -322 64
rect -305 62 -299 64
rect -329 60 -326 62
rect -324 60 -322 62
rect -329 51 -322 60
rect -314 57 -309 62
rect -316 55 -309 57
rect -316 53 -314 55
rect -312 53 -309 55
rect -349 44 -343 51
rect -316 48 -309 53
rect -316 46 -314 48
rect -312 46 -309 48
rect -316 44 -309 46
rect -307 60 -299 62
rect -307 58 -304 60
rect -302 58 -299 60
rect -307 51 -299 58
rect -297 62 -289 64
rect -297 60 -294 62
rect -292 60 -289 62
rect -297 55 -289 60
rect -297 53 -294 55
rect -292 53 -289 55
rect -297 51 -289 53
rect -287 62 -280 64
rect -261 62 -255 64
rect -287 60 -284 62
rect -282 60 -280 62
rect -287 51 -280 60
rect -270 57 -265 62
rect -272 55 -265 57
rect -272 53 -270 55
rect -268 53 -265 55
rect -307 44 -301 51
rect -272 48 -265 53
rect -272 46 -270 48
rect -268 46 -265 48
rect -272 44 -265 46
rect -263 60 -255 62
rect -263 58 -260 60
rect -258 58 -255 60
rect -263 51 -255 58
rect -253 62 -245 64
rect -253 60 -250 62
rect -248 60 -245 62
rect -253 55 -245 60
rect -253 53 -250 55
rect -248 53 -245 55
rect -253 51 -245 53
rect -243 62 -236 64
rect -192 62 -186 64
rect -243 60 -240 62
rect -238 60 -236 62
rect -243 51 -236 60
rect -201 57 -196 62
rect -203 55 -196 57
rect -203 53 -201 55
rect -199 53 -196 55
rect -263 44 -257 51
rect -203 48 -196 53
rect -203 46 -201 48
rect -199 46 -196 48
rect -203 44 -196 46
rect -194 60 -186 62
rect -194 58 -191 60
rect -189 58 -186 60
rect -194 51 -186 58
rect -184 62 -176 64
rect -184 60 -181 62
rect -179 60 -176 62
rect -184 55 -176 60
rect -184 53 -181 55
rect -179 53 -176 55
rect -184 51 -176 53
rect -174 62 -167 64
rect -148 62 -142 64
rect -174 60 -171 62
rect -169 60 -167 62
rect -174 51 -167 60
rect -157 57 -152 62
rect -159 55 -152 57
rect -159 53 -157 55
rect -155 53 -152 55
rect -194 44 -188 51
rect -159 48 -152 53
rect -159 46 -157 48
rect -155 46 -152 48
rect -159 44 -152 46
rect -150 60 -142 62
rect -150 58 -147 60
rect -145 58 -142 60
rect -150 51 -142 58
rect -140 62 -132 64
rect -140 60 -137 62
rect -135 60 -132 62
rect -140 55 -132 60
rect -140 53 -137 55
rect -135 53 -132 55
rect -140 51 -132 53
rect -130 62 -123 64
rect -106 62 -100 64
rect -130 60 -127 62
rect -125 60 -123 62
rect -130 51 -123 60
rect -115 57 -110 62
rect -117 55 -110 57
rect -117 53 -115 55
rect -113 53 -110 55
rect -150 44 -144 51
rect -117 48 -110 53
rect -117 46 -115 48
rect -113 46 -110 48
rect -117 44 -110 46
rect -108 60 -100 62
rect -108 58 -105 60
rect -103 58 -100 60
rect -108 51 -100 58
rect -98 62 -90 64
rect -98 60 -95 62
rect -93 60 -90 62
rect -98 55 -90 60
rect -98 53 -95 55
rect -93 53 -90 55
rect -98 51 -90 53
rect -88 62 -81 64
rect -65 62 -59 64
rect -88 60 -85 62
rect -83 60 -81 62
rect -88 51 -81 60
rect -74 57 -69 62
rect -76 55 -69 57
rect -76 53 -74 55
rect -72 53 -69 55
rect -108 44 -102 51
rect -76 48 -69 53
rect -76 46 -74 48
rect -72 46 -69 48
rect -76 44 -69 46
rect -67 60 -59 62
rect -67 58 -64 60
rect -62 58 -59 60
rect -67 51 -59 58
rect -57 62 -49 64
rect -57 60 -54 62
rect -52 60 -49 62
rect -57 55 -49 60
rect -57 53 -54 55
rect -52 53 -49 55
rect -57 51 -49 53
rect -47 62 -40 64
rect -22 62 -16 64
rect -47 60 -44 62
rect -42 60 -40 62
rect -47 51 -40 60
rect -31 57 -26 62
rect -33 55 -26 57
rect -33 53 -31 55
rect -29 53 -26 55
rect -67 44 -61 51
rect -33 48 -26 53
rect -33 46 -31 48
rect -29 46 -26 48
rect -33 44 -26 46
rect -24 60 -16 62
rect -24 58 -21 60
rect -19 58 -16 60
rect -24 51 -16 58
rect -14 62 -6 64
rect -14 60 -11 62
rect -9 60 -6 62
rect -14 55 -6 60
rect -14 53 -11 55
rect -9 53 -6 55
rect -14 51 -6 53
rect -4 62 3 64
rect 18 62 24 64
rect -4 60 -1 62
rect 1 60 3 62
rect -4 51 3 60
rect 9 57 14 62
rect 7 55 14 57
rect 7 53 9 55
rect 11 53 14 55
rect -24 44 -18 51
rect 7 48 14 53
rect 7 46 9 48
rect 11 46 14 48
rect 7 44 14 46
rect 16 60 24 62
rect 16 58 19 60
rect 21 58 24 60
rect 16 51 24 58
rect 26 62 34 64
rect 26 60 29 62
rect 31 60 34 62
rect 26 55 34 60
rect 26 53 29 55
rect 31 53 34 55
rect 26 51 34 53
rect 36 62 43 64
rect 61 62 67 64
rect 36 60 39 62
rect 41 60 43 62
rect 36 51 43 60
rect 52 57 57 62
rect 50 55 57 57
rect 50 53 52 55
rect 54 53 57 55
rect 16 44 22 51
rect 50 48 57 53
rect 50 46 52 48
rect 54 46 57 48
rect 50 44 57 46
rect 59 60 67 62
rect 59 58 62 60
rect 64 58 67 60
rect 59 51 67 58
rect 69 62 77 64
rect 69 60 72 62
rect 74 60 77 62
rect 69 55 77 60
rect 69 53 72 55
rect 74 53 77 55
rect 69 51 77 53
rect 79 62 86 64
rect 79 60 82 62
rect 84 60 86 62
rect 79 51 86 60
rect 59 44 65 51
rect -572 -34 -565 -32
rect -572 -36 -570 -34
rect -568 -36 -565 -34
rect -572 -41 -565 -36
rect -572 -43 -570 -41
rect -568 -43 -565 -41
rect -572 -45 -565 -43
rect -570 -60 -565 -45
rect -563 -49 -555 -32
rect -563 -51 -560 -49
rect -558 -51 -555 -49
rect -563 -56 -555 -51
rect -563 -58 -560 -56
rect -558 -58 -555 -56
rect -563 -60 -555 -58
rect -553 -41 -545 -32
rect -553 -43 -550 -41
rect -548 -43 -545 -41
rect -553 -48 -545 -43
rect -553 -50 -550 -48
rect -548 -50 -545 -48
rect -553 -60 -545 -50
rect -543 -49 -527 -32
rect -543 -51 -538 -49
rect -536 -51 -527 -49
rect -543 -56 -527 -51
rect -543 -58 -538 -56
rect -536 -57 -527 -56
rect -525 -57 -520 -32
rect -518 -35 -513 -32
rect -481 -34 -474 -32
rect -518 -37 -510 -35
rect -518 -39 -515 -37
rect -513 -39 -510 -37
rect -518 -48 -510 -39
rect -508 -48 -497 -35
rect -518 -57 -513 -48
rect -506 -56 -497 -48
rect -536 -58 -529 -57
rect -543 -60 -529 -58
rect -506 -58 -503 -56
rect -501 -58 -497 -56
rect -506 -60 -497 -58
rect -495 -37 -488 -35
rect -495 -39 -492 -37
rect -490 -39 -488 -37
rect -495 -44 -488 -39
rect -495 -46 -492 -44
rect -490 -46 -488 -44
rect -481 -36 -479 -34
rect -477 -36 -474 -34
rect -481 -41 -474 -36
rect -481 -43 -479 -41
rect -477 -43 -474 -41
rect -481 -45 -474 -43
rect -495 -48 -488 -46
rect -495 -60 -490 -48
rect -479 -50 -474 -45
rect -472 -49 -463 -32
rect -452 -40 -447 -32
rect -472 -50 -468 -49
rect -470 -51 -468 -50
rect -466 -51 -463 -49
rect -470 -53 -463 -51
rect -454 -42 -447 -40
rect -454 -44 -452 -42
rect -450 -44 -447 -42
rect -454 -49 -447 -44
rect -454 -51 -452 -49
rect -450 -51 -447 -49
rect -454 -53 -447 -51
rect -452 -59 -447 -53
rect -445 -48 -437 -32
rect -445 -50 -442 -48
rect -440 -50 -437 -48
rect -445 -55 -437 -50
rect -445 -57 -442 -55
rect -440 -57 -437 -55
rect -445 -59 -437 -57
rect -435 -59 -430 -32
rect -428 -34 -420 -32
rect -428 -36 -425 -34
rect -423 -36 -420 -34
rect -428 -41 -420 -36
rect -428 -43 -425 -41
rect -423 -43 -420 -41
rect -428 -59 -420 -43
rect -418 -50 -410 -32
rect -418 -52 -415 -50
rect -413 -52 -410 -50
rect -418 -59 -410 -52
rect -408 -47 -401 -32
rect -390 -47 -385 -32
rect -408 -49 -405 -47
rect -403 -49 -401 -47
rect -408 -55 -401 -49
rect -392 -49 -385 -47
rect -392 -51 -390 -49
rect -388 -51 -385 -49
rect -392 -53 -385 -51
rect -408 -57 -405 -55
rect -403 -57 -401 -55
rect -408 -59 -401 -57
rect -390 -60 -385 -53
rect -383 -41 -375 -32
rect -383 -43 -380 -41
rect -378 -43 -375 -41
rect -383 -60 -375 -43
rect -373 -34 -365 -32
rect -373 -36 -370 -34
rect -368 -36 -365 -34
rect -373 -41 -365 -36
rect -373 -43 -370 -41
rect -368 -43 -365 -41
rect -373 -60 -365 -43
rect -363 -46 -357 -32
rect -363 -56 -355 -46
rect -363 -58 -360 -56
rect -358 -58 -355 -56
rect -363 -60 -355 -58
rect -353 -49 -345 -46
rect -353 -51 -350 -49
rect -348 -51 -345 -49
rect -353 -60 -345 -51
rect -343 -49 -336 -46
rect -330 -47 -325 -32
rect -343 -51 -340 -49
rect -338 -51 -336 -49
rect -343 -56 -336 -51
rect -332 -49 -325 -47
rect -332 -51 -330 -49
rect -328 -51 -325 -49
rect -332 -53 -325 -51
rect -343 -58 -340 -56
rect -338 -58 -336 -56
rect -343 -60 -336 -58
rect -330 -60 -325 -53
rect -323 -41 -315 -32
rect -323 -43 -320 -41
rect -318 -43 -315 -41
rect -323 -60 -315 -43
rect -313 -34 -305 -32
rect -313 -36 -310 -34
rect -308 -36 -305 -34
rect -313 -41 -305 -36
rect -313 -43 -310 -41
rect -308 -43 -305 -41
rect -313 -60 -305 -43
rect -303 -39 -296 -32
rect -263 -34 -256 -32
rect -263 -36 -261 -34
rect -259 -36 -256 -34
rect -303 -53 -294 -39
rect -292 -41 -284 -39
rect -292 -43 -289 -41
rect -287 -43 -284 -41
rect -292 -53 -284 -43
rect -282 -49 -274 -39
rect -263 -41 -256 -36
rect -263 -43 -261 -41
rect -259 -43 -256 -41
rect -263 -45 -256 -43
rect -282 -51 -279 -49
rect -277 -51 -274 -49
rect -261 -50 -256 -45
rect -254 -49 -245 -32
rect -234 -40 -229 -32
rect -254 -50 -250 -49
rect -282 -53 -274 -51
rect -303 -56 -296 -53
rect -303 -58 -300 -56
rect -298 -58 -296 -56
rect -252 -51 -250 -50
rect -248 -51 -245 -49
rect -252 -53 -245 -51
rect -236 -42 -229 -40
rect -236 -44 -234 -42
rect -232 -44 -229 -42
rect -236 -49 -229 -44
rect -236 -51 -234 -49
rect -232 -51 -229 -49
rect -236 -53 -229 -51
rect -303 -60 -296 -58
rect -234 -59 -229 -53
rect -227 -48 -219 -32
rect -227 -50 -224 -48
rect -222 -50 -219 -48
rect -227 -55 -219 -50
rect -227 -57 -224 -55
rect -222 -57 -219 -55
rect -227 -59 -219 -57
rect -217 -59 -212 -32
rect -210 -34 -202 -32
rect -210 -36 -207 -34
rect -205 -36 -202 -34
rect -210 -41 -202 -36
rect -210 -43 -207 -41
rect -205 -43 -202 -41
rect -210 -59 -202 -43
rect -200 -50 -192 -32
rect -200 -52 -197 -50
rect -195 -52 -192 -50
rect -200 -59 -192 -52
rect -190 -47 -183 -32
rect -172 -47 -167 -32
rect -190 -49 -187 -47
rect -185 -49 -183 -47
rect -190 -55 -183 -49
rect -174 -49 -167 -47
rect -174 -51 -172 -49
rect -170 -51 -167 -49
rect -174 -53 -167 -51
rect -190 -57 -187 -55
rect -185 -57 -183 -55
rect -190 -59 -183 -57
rect -172 -60 -167 -53
rect -165 -41 -157 -32
rect -165 -43 -162 -41
rect -160 -43 -157 -41
rect -165 -60 -157 -43
rect -155 -34 -147 -32
rect -155 -36 -152 -34
rect -150 -36 -147 -34
rect -155 -41 -147 -36
rect -155 -43 -152 -41
rect -150 -43 -147 -41
rect -155 -60 -147 -43
rect -145 -46 -139 -32
rect -145 -56 -137 -46
rect -145 -58 -142 -56
rect -140 -58 -137 -56
rect -145 -60 -137 -58
rect -135 -49 -127 -46
rect -135 -51 -132 -49
rect -130 -51 -127 -49
rect -135 -60 -127 -51
rect -125 -49 -118 -46
rect -112 -47 -107 -32
rect -125 -51 -122 -49
rect -120 -51 -118 -49
rect -125 -56 -118 -51
rect -114 -49 -107 -47
rect -114 -51 -112 -49
rect -110 -51 -107 -49
rect -114 -53 -107 -51
rect -125 -58 -122 -56
rect -120 -58 -118 -56
rect -125 -60 -118 -58
rect -112 -60 -107 -53
rect -105 -41 -97 -32
rect -105 -43 -102 -41
rect -100 -43 -97 -41
rect -105 -60 -97 -43
rect -95 -34 -87 -32
rect -95 -36 -92 -34
rect -90 -36 -87 -34
rect -95 -41 -87 -36
rect -95 -43 -92 -41
rect -90 -43 -87 -41
rect -95 -60 -87 -43
rect -85 -39 -78 -32
rect -34 -34 -27 -32
rect -34 -36 -32 -34
rect -30 -36 -27 -34
rect -85 -53 -76 -39
rect -74 -41 -66 -39
rect -74 -43 -71 -41
rect -69 -43 -66 -41
rect -74 -53 -66 -43
rect -64 -49 -56 -39
rect -34 -41 -27 -36
rect -34 -43 -32 -41
rect -30 -43 -27 -41
rect -34 -45 -27 -43
rect -64 -51 -61 -49
rect -59 -51 -56 -49
rect -64 -53 -56 -51
rect -85 -56 -78 -53
rect -85 -58 -82 -56
rect -80 -58 -78 -56
rect -85 -60 -78 -58
rect -32 -60 -27 -45
rect -25 -49 -17 -32
rect -25 -51 -22 -49
rect -20 -51 -17 -49
rect -25 -56 -17 -51
rect -25 -58 -22 -56
rect -20 -58 -17 -56
rect -25 -60 -17 -58
rect -15 -41 -7 -32
rect -15 -43 -12 -41
rect -10 -43 -7 -41
rect -15 -48 -7 -43
rect -15 -50 -12 -48
rect -10 -50 -7 -48
rect -15 -60 -7 -50
rect -5 -49 11 -32
rect -5 -51 0 -49
rect 2 -51 11 -49
rect -5 -56 11 -51
rect -5 -58 0 -56
rect 2 -57 11 -56
rect 13 -57 18 -32
rect 20 -35 25 -32
rect 20 -37 28 -35
rect 20 -39 23 -37
rect 25 -39 28 -37
rect 20 -48 28 -39
rect 30 -48 41 -35
rect 20 -57 25 -48
rect 32 -56 41 -48
rect 2 -58 9 -57
rect -5 -60 9 -58
rect 32 -58 35 -56
rect 37 -58 41 -56
rect 32 -60 41 -58
rect 43 -37 50 -35
rect 43 -39 46 -37
rect 48 -39 50 -37
rect 43 -44 50 -39
rect 43 -46 46 -44
rect 48 -46 50 -44
rect 43 -48 50 -46
rect 43 -60 48 -48
rect -488 -79 -483 -73
rect -506 -81 -499 -79
rect -506 -82 -504 -81
rect -515 -87 -510 -82
rect -517 -89 -510 -87
rect -517 -91 -515 -89
rect -513 -91 -510 -89
rect -517 -96 -510 -91
rect -517 -98 -515 -96
rect -513 -98 -510 -96
rect -517 -100 -510 -98
rect -508 -83 -504 -82
rect -502 -83 -499 -81
rect -508 -100 -499 -83
rect -490 -81 -483 -79
rect -490 -83 -488 -81
rect -486 -83 -483 -81
rect -490 -88 -483 -83
rect -490 -90 -488 -88
rect -486 -90 -483 -88
rect -490 -92 -483 -90
rect -488 -100 -483 -92
rect -481 -75 -473 -73
rect -481 -77 -478 -75
rect -476 -77 -473 -75
rect -481 -82 -473 -77
rect -481 -84 -478 -82
rect -476 -84 -473 -82
rect -481 -100 -473 -84
rect -471 -100 -466 -73
rect -464 -89 -456 -73
rect -464 -91 -461 -89
rect -459 -91 -456 -89
rect -464 -96 -456 -91
rect -464 -98 -461 -96
rect -459 -98 -456 -96
rect -464 -100 -456 -98
rect -454 -80 -446 -73
rect -454 -82 -451 -80
rect -449 -82 -446 -80
rect -454 -100 -446 -82
rect -444 -75 -437 -73
rect -444 -77 -441 -75
rect -439 -77 -437 -75
rect -444 -83 -437 -77
rect -426 -79 -421 -72
rect -444 -85 -441 -83
rect -439 -85 -437 -83
rect -428 -81 -421 -79
rect -428 -83 -426 -81
rect -424 -83 -421 -81
rect -428 -85 -421 -83
rect -444 -100 -437 -85
rect -426 -100 -421 -85
rect -419 -89 -411 -72
rect -419 -91 -416 -89
rect -414 -91 -411 -89
rect -419 -100 -411 -91
rect -409 -89 -401 -72
rect -409 -91 -406 -89
rect -404 -91 -401 -89
rect -409 -96 -401 -91
rect -409 -98 -406 -96
rect -404 -98 -401 -96
rect -409 -100 -401 -98
rect -399 -74 -391 -72
rect -399 -76 -396 -74
rect -394 -76 -391 -74
rect -399 -86 -391 -76
rect -389 -81 -381 -72
rect -389 -83 -386 -81
rect -384 -83 -381 -81
rect -389 -86 -381 -83
rect -379 -74 -372 -72
rect -379 -76 -376 -74
rect -374 -76 -372 -74
rect -379 -81 -372 -76
rect -366 -79 -361 -72
rect -379 -83 -376 -81
rect -374 -83 -372 -81
rect -379 -86 -372 -83
rect -368 -81 -361 -79
rect -368 -83 -366 -81
rect -364 -83 -361 -81
rect -368 -85 -361 -83
rect -399 -100 -393 -86
rect -366 -100 -361 -85
rect -359 -89 -351 -72
rect -359 -91 -356 -89
rect -354 -91 -351 -89
rect -359 -100 -351 -91
rect -349 -89 -341 -72
rect -349 -91 -346 -89
rect -344 -91 -341 -89
rect -349 -96 -341 -91
rect -349 -98 -346 -96
rect -344 -98 -341 -96
rect -349 -100 -341 -98
rect -339 -74 -332 -72
rect -339 -76 -336 -74
rect -334 -76 -332 -74
rect -339 -79 -332 -76
rect -339 -93 -330 -79
rect -328 -89 -320 -79
rect -328 -91 -325 -89
rect -323 -91 -320 -89
rect -328 -93 -320 -91
rect -318 -81 -310 -79
rect -318 -83 -315 -81
rect -313 -83 -310 -81
rect -268 -79 -263 -73
rect -286 -81 -279 -79
rect -286 -82 -284 -81
rect -318 -93 -310 -83
rect -295 -87 -290 -82
rect -297 -89 -290 -87
rect -297 -91 -295 -89
rect -293 -91 -290 -89
rect -339 -100 -332 -93
rect -297 -96 -290 -91
rect -297 -98 -295 -96
rect -293 -98 -290 -96
rect -297 -100 -290 -98
rect -288 -83 -284 -82
rect -282 -83 -279 -81
rect -288 -100 -279 -83
rect -270 -81 -263 -79
rect -270 -83 -268 -81
rect -266 -83 -263 -81
rect -270 -88 -263 -83
rect -270 -90 -268 -88
rect -266 -90 -263 -88
rect -270 -92 -263 -90
rect -268 -100 -263 -92
rect -261 -75 -253 -73
rect -261 -77 -258 -75
rect -256 -77 -253 -75
rect -261 -82 -253 -77
rect -261 -84 -258 -82
rect -256 -84 -253 -82
rect -261 -100 -253 -84
rect -251 -100 -246 -73
rect -244 -89 -236 -73
rect -244 -91 -241 -89
rect -239 -91 -236 -89
rect -244 -96 -236 -91
rect -244 -98 -241 -96
rect -239 -98 -236 -96
rect -244 -100 -236 -98
rect -234 -80 -226 -73
rect -234 -82 -231 -80
rect -229 -82 -226 -80
rect -234 -100 -226 -82
rect -224 -75 -217 -73
rect -224 -77 -221 -75
rect -219 -77 -217 -75
rect -224 -83 -217 -77
rect -206 -79 -201 -72
rect -224 -85 -221 -83
rect -219 -85 -217 -83
rect -208 -81 -201 -79
rect -208 -83 -206 -81
rect -204 -83 -201 -81
rect -208 -85 -201 -83
rect -224 -100 -217 -85
rect -206 -100 -201 -85
rect -199 -89 -191 -72
rect -199 -91 -196 -89
rect -194 -91 -191 -89
rect -199 -100 -191 -91
rect -189 -89 -181 -72
rect -189 -91 -186 -89
rect -184 -91 -181 -89
rect -189 -96 -181 -91
rect -189 -98 -186 -96
rect -184 -98 -181 -96
rect -189 -100 -181 -98
rect -179 -74 -171 -72
rect -179 -76 -176 -74
rect -174 -76 -171 -74
rect -179 -86 -171 -76
rect -169 -81 -161 -72
rect -169 -83 -166 -81
rect -164 -83 -161 -81
rect -169 -86 -161 -83
rect -159 -74 -152 -72
rect -159 -76 -156 -74
rect -154 -76 -152 -74
rect -159 -81 -152 -76
rect -146 -79 -141 -72
rect -159 -83 -156 -81
rect -154 -83 -152 -81
rect -159 -86 -152 -83
rect -148 -81 -141 -79
rect -148 -83 -146 -81
rect -144 -83 -141 -81
rect -148 -85 -141 -83
rect -179 -100 -173 -86
rect -146 -100 -141 -85
rect -139 -89 -131 -72
rect -139 -91 -136 -89
rect -134 -91 -131 -89
rect -139 -100 -131 -91
rect -129 -89 -121 -72
rect -129 -91 -126 -89
rect -124 -91 -121 -89
rect -129 -96 -121 -91
rect -129 -98 -126 -96
rect -124 -98 -121 -96
rect -129 -100 -121 -98
rect -119 -74 -112 -72
rect -119 -76 -116 -74
rect -114 -76 -112 -74
rect -119 -79 -112 -76
rect -119 -93 -110 -79
rect -108 -89 -100 -79
rect -108 -91 -105 -89
rect -103 -91 -100 -89
rect -108 -93 -100 -91
rect -98 -81 -90 -79
rect -98 -83 -95 -81
rect -93 -83 -90 -81
rect -98 -93 -90 -83
rect -73 -87 -68 -72
rect -75 -89 -68 -87
rect -75 -91 -73 -89
rect -71 -91 -68 -89
rect -119 -100 -112 -93
rect -75 -96 -68 -91
rect -75 -98 -73 -96
rect -71 -98 -68 -96
rect -75 -100 -68 -98
rect -66 -74 -58 -72
rect -66 -76 -63 -74
rect -61 -76 -58 -74
rect -66 -81 -58 -76
rect -66 -83 -63 -81
rect -61 -83 -58 -81
rect -66 -100 -58 -83
rect -56 -82 -48 -72
rect -56 -84 -53 -82
rect -51 -84 -48 -82
rect -56 -89 -48 -84
rect -56 -91 -53 -89
rect -51 -91 -48 -89
rect -56 -100 -48 -91
rect -46 -74 -32 -72
rect -46 -76 -41 -74
rect -39 -75 -32 -74
rect -9 -74 0 -72
rect -39 -76 -30 -75
rect -46 -81 -30 -76
rect -46 -83 -41 -81
rect -39 -83 -30 -81
rect -46 -100 -30 -83
rect -28 -100 -23 -75
rect -21 -84 -16 -75
rect -9 -76 -6 -74
rect -4 -76 0 -74
rect -9 -84 0 -76
rect -21 -93 -13 -84
rect -21 -95 -18 -93
rect -16 -95 -13 -93
rect -21 -97 -13 -95
rect -11 -97 0 -84
rect 2 -84 7 -72
rect 2 -86 9 -84
rect 2 -88 5 -86
rect 7 -88 9 -86
rect 2 -93 9 -88
rect 2 -95 5 -93
rect 7 -95 9 -93
rect 2 -97 9 -95
rect -21 -100 -16 -97
<< alu1 >>
rect -549 72 90 77
rect -549 70 -542 72
rect -540 70 -502 72
rect -500 70 -459 72
rect -457 70 -355 72
rect -353 70 -313 72
rect -311 70 -269 72
rect -267 70 -200 72
rect -198 70 -156 72
rect -154 70 -114 72
rect -112 70 -73 72
rect -71 70 -30 72
rect -28 70 10 72
rect 12 70 53 72
rect 55 70 90 72
rect -549 69 90 70
rect -545 55 -540 57
rect -545 53 -543 55
rect -541 53 -540 55
rect -545 48 -540 53
rect -545 46 -543 48
rect -541 46 -540 48
rect -545 44 -540 46
rect -513 55 -509 56
rect -513 53 -512 55
rect -510 53 -509 55
rect -545 24 -541 44
rect -513 47 -509 53
rect -522 46 -509 47
rect -522 44 -516 46
rect -514 44 -509 46
rect -522 43 -509 44
rect -505 55 -500 57
rect -505 53 -503 55
rect -501 53 -500 55
rect -505 48 -500 53
rect -505 46 -503 48
rect -501 46 -500 48
rect -505 44 -500 46
rect -473 55 -469 56
rect -473 53 -472 55
rect -470 53 -469 55
rect -530 38 -516 39
rect -530 36 -526 38
rect -524 37 -516 38
rect -524 36 -520 37
rect -530 35 -520 36
rect -518 35 -516 37
rect -545 22 -543 24
rect -541 22 -533 24
rect -545 21 -533 22
rect -545 19 -539 21
rect -537 19 -533 21
rect -521 26 -516 35
rect -505 24 -501 44
rect -473 47 -469 53
rect -482 46 -469 47
rect -482 44 -476 46
rect -474 44 -469 46
rect -482 43 -469 44
rect -462 55 -457 57
rect -462 53 -460 55
rect -458 53 -457 55
rect -462 48 -457 53
rect -462 46 -460 48
rect -458 46 -457 48
rect -462 44 -457 46
rect -430 50 -426 56
rect -490 38 -476 39
rect -490 36 -486 38
rect -484 36 -480 38
rect -478 36 -476 38
rect -490 35 -476 36
rect -505 22 -503 24
rect -501 22 -493 24
rect -505 21 -493 22
rect -505 19 -503 21
rect -501 19 -493 21
rect -481 26 -476 35
rect -462 24 -458 44
rect -430 48 -429 50
rect -427 48 -426 50
rect -430 47 -426 48
rect -439 46 -426 47
rect -439 44 -433 46
rect -431 44 -426 46
rect -439 43 -426 44
rect -358 55 -353 57
rect -358 53 -356 55
rect -354 53 -353 55
rect -358 48 -353 53
rect -358 46 -356 48
rect -354 46 -353 48
rect -358 44 -353 46
rect -326 50 -322 56
rect -447 38 -433 39
rect -447 36 -443 38
rect -441 36 -433 38
rect -447 35 -433 36
rect -462 22 -460 24
rect -458 22 -450 24
rect -462 21 -450 22
rect -462 19 -460 21
rect -458 19 -450 21
rect -438 29 -433 35
rect -438 27 -436 29
rect -434 27 -433 29
rect -438 26 -433 27
rect -358 24 -354 44
rect -326 48 -325 50
rect -323 48 -322 50
rect -326 47 -322 48
rect -335 46 -322 47
rect -335 44 -329 46
rect -327 44 -322 46
rect -335 43 -322 44
rect -316 55 -311 57
rect -316 53 -314 55
rect -312 53 -311 55
rect -316 48 -311 53
rect -316 46 -314 48
rect -312 46 -311 48
rect -316 44 -311 46
rect -284 55 -280 56
rect -284 53 -283 55
rect -281 53 -280 55
rect -343 38 -329 39
rect -343 36 -339 38
rect -337 36 -329 38
rect -343 35 -329 36
rect -358 22 -356 24
rect -354 22 -346 24
rect -358 21 -346 22
rect -358 19 -353 21
rect -351 19 -346 21
rect -334 30 -329 35
rect -334 28 -333 30
rect -331 28 -329 30
rect -334 26 -329 28
rect -316 24 -312 44
rect -284 47 -280 53
rect -293 46 -280 47
rect -293 44 -287 46
rect -285 44 -280 46
rect -293 43 -280 44
rect -272 55 -267 57
rect -272 53 -270 55
rect -268 53 -267 55
rect -272 48 -267 53
rect -272 46 -270 48
rect -268 46 -267 48
rect -272 44 -267 46
rect -240 55 -236 56
rect -240 53 -239 55
rect -237 53 -236 55
rect -301 38 -287 39
rect -301 36 -297 38
rect -295 36 -291 38
rect -289 36 -287 38
rect -301 35 -287 36
rect -316 22 -314 24
rect -312 22 -304 24
rect -316 21 -304 22
rect -316 19 -315 21
rect -313 19 -304 21
rect -292 26 -287 35
rect -272 30 -268 44
rect -272 28 -271 30
rect -269 28 -268 30
rect -272 24 -268 28
rect -240 47 -236 53
rect -249 46 -236 47
rect -249 44 -243 46
rect -241 44 -236 46
rect -249 43 -236 44
rect -203 55 -198 57
rect -203 53 -201 55
rect -199 53 -198 55
rect -203 48 -198 53
rect -203 46 -201 48
rect -199 46 -198 48
rect -203 44 -198 46
rect -171 55 -167 56
rect -171 53 -170 55
rect -168 53 -167 55
rect -257 38 -243 39
rect -257 36 -253 38
rect -251 36 -243 38
rect -257 35 -243 36
rect -272 22 -270 24
rect -268 22 -260 24
rect -545 18 -533 19
rect -505 18 -493 19
rect -462 18 -450 19
rect -358 18 -346 19
rect -316 18 -304 19
rect -272 18 -260 22
rect -248 30 -243 35
rect -248 28 -247 30
rect -245 28 -243 30
rect -248 26 -243 28
rect -203 24 -199 44
rect -171 47 -167 53
rect -180 46 -167 47
rect -180 44 -174 46
rect -172 44 -167 46
rect -180 43 -167 44
rect -159 55 -154 57
rect -159 53 -157 55
rect -155 53 -154 55
rect -159 48 -154 53
rect -159 46 -157 48
rect -155 46 -154 48
rect -159 44 -154 46
rect -127 55 -123 56
rect -127 53 -126 55
rect -124 53 -123 55
rect -188 38 -174 39
rect -188 36 -184 38
rect -182 36 -174 38
rect -188 35 -174 36
rect -203 22 -201 24
rect -199 22 -191 24
rect -203 21 -191 22
rect -203 19 -199 21
rect -197 19 -191 21
rect -179 30 -174 35
rect -179 28 -178 30
rect -176 28 -174 30
rect -179 26 -174 28
rect -159 24 -155 44
rect -127 47 -123 53
rect -136 46 -123 47
rect -136 44 -130 46
rect -128 44 -123 46
rect -136 43 -123 44
rect -117 55 -112 57
rect -117 53 -115 55
rect -113 53 -112 55
rect -117 48 -112 53
rect -117 46 -115 48
rect -113 46 -112 48
rect -117 44 -112 46
rect -85 50 -81 56
rect -144 38 -130 39
rect -144 36 -140 38
rect -138 36 -130 38
rect -144 35 -130 36
rect -159 22 -157 24
rect -155 22 -147 24
rect -159 20 -150 22
rect -148 20 -147 22
rect -203 18 -191 19
rect -159 18 -147 20
rect -135 30 -130 35
rect -135 28 -134 30
rect -132 28 -130 30
rect -135 26 -130 28
rect -117 24 -113 44
rect -85 48 -84 50
rect -82 48 -81 50
rect -85 47 -81 48
rect -94 46 -81 47
rect -94 44 -88 46
rect -86 44 -81 46
rect -94 43 -81 44
rect -76 55 -71 57
rect -76 53 -74 55
rect -72 53 -71 55
rect -76 48 -71 53
rect -76 46 -74 48
rect -72 46 -71 48
rect -76 44 -71 46
rect -44 54 -40 56
rect -44 52 -43 54
rect -41 52 -40 54
rect -102 38 -88 39
rect -102 36 -98 38
rect -96 36 -92 38
rect -90 36 -88 38
rect -102 35 -88 36
rect -117 22 -115 24
rect -113 22 -105 24
rect -117 21 -105 22
rect -117 19 -116 21
rect -114 19 -105 21
rect -93 26 -88 35
rect -76 24 -72 44
rect -44 47 -40 52
rect -53 46 -40 47
rect -53 44 -47 46
rect -45 44 -40 46
rect -53 43 -40 44
rect -33 55 -28 57
rect -33 53 -31 55
rect -29 53 -28 55
rect -33 48 -28 53
rect -33 46 -31 48
rect -29 46 -28 48
rect -33 44 -28 46
rect -1 55 3 56
rect -1 53 0 55
rect 2 53 3 55
rect -61 38 -47 39
rect -61 36 -57 38
rect -55 36 -47 38
rect -61 35 -47 36
rect -76 22 -74 24
rect -72 22 -64 24
rect -76 21 -64 22
rect -76 19 -68 21
rect -66 19 -64 21
rect -52 30 -47 35
rect -52 28 -51 30
rect -49 28 -47 30
rect -52 26 -47 28
rect -33 24 -29 44
rect -1 47 3 53
rect -10 46 3 47
rect -10 44 -4 46
rect -2 44 3 46
rect -10 43 3 44
rect 7 55 12 57
rect 7 53 9 55
rect 11 53 12 55
rect 7 48 12 53
rect 7 46 9 48
rect 11 46 12 48
rect 7 44 12 46
rect 39 50 43 56
rect -18 38 -4 39
rect -18 36 -14 38
rect -12 36 -8 38
rect -6 36 -4 38
rect -18 35 -4 36
rect -33 22 -31 24
rect -29 22 -21 24
rect -33 21 -21 22
rect -33 19 -25 21
rect -23 19 -21 21
rect -9 26 -4 35
rect 7 24 11 44
rect 39 48 40 50
rect 42 48 43 50
rect 39 47 43 48
rect 30 46 43 47
rect 30 44 36 46
rect 38 44 43 46
rect 30 43 43 44
rect 50 55 55 57
rect 50 53 52 55
rect 54 53 55 55
rect 50 48 55 53
rect 50 46 52 48
rect 54 46 55 48
rect 50 44 55 46
rect 82 55 86 56
rect 82 53 83 55
rect 85 53 86 55
rect 22 38 36 39
rect 22 36 26 38
rect 28 36 36 38
rect 22 35 36 36
rect 7 22 9 24
rect 11 22 19 24
rect 7 21 19 22
rect 7 19 15 21
rect 17 19 19 21
rect 31 29 36 35
rect 31 27 33 29
rect 35 27 36 29
rect 31 26 36 27
rect 50 24 54 44
rect 82 47 86 53
rect 73 46 86 47
rect 73 44 79 46
rect 81 44 86 46
rect 73 43 86 44
rect 65 38 79 39
rect 65 36 69 38
rect 71 36 79 38
rect 65 35 79 36
rect 50 22 52 24
rect 54 22 62 24
rect -117 18 -105 19
rect -76 18 -64 19
rect -33 18 -21 19
rect 7 18 19 19
rect 50 18 62 22
rect 74 29 79 35
rect 74 27 76 29
rect 78 27 79 29
rect 74 26 79 27
rect -549 12 90 13
rect -549 10 -542 12
rect -540 10 -532 12
rect -530 10 -502 12
rect -500 10 -492 12
rect -490 10 -459 12
rect -457 10 -449 12
rect -447 10 -355 12
rect -353 10 -345 12
rect -343 10 -313 12
rect -311 10 -303 12
rect -301 10 -269 12
rect -267 10 -259 12
rect -257 10 -200 12
rect -198 10 -190 12
rect -188 10 -156 12
rect -154 10 -146 12
rect -144 10 -114 12
rect -112 10 -104 12
rect -102 10 -73 12
rect -71 10 -63 12
rect -61 10 -30 12
rect -28 10 -20 12
rect -18 10 10 12
rect 12 10 20 12
rect 22 10 53 12
rect 55 10 63 12
rect 65 10 90 12
rect -549 6 90 10
rect -584 5 90 6
rect -584 1 54 5
rect -584 -1 -478 1
rect -476 -1 -466 1
rect -464 -1 -444 1
rect -442 -1 -390 1
rect -388 -1 -328 1
rect -326 -1 -273 1
rect -271 -1 -260 1
rect -258 -1 -248 1
rect -246 -1 -226 1
rect -224 -1 -172 1
rect -170 -1 -110 1
rect -108 -1 -55 1
rect -53 -1 54 1
rect -584 -2 54 -1
rect -573 -9 -551 -8
rect -573 -11 -570 -9
rect -568 -11 -551 -9
rect -573 -12 -551 -11
rect -493 -9 -488 -7
rect -493 -11 -492 -9
rect -490 -11 -488 -9
rect -573 -32 -569 -12
rect -540 -17 -536 -15
rect -540 -19 -539 -17
rect -537 -19 -536 -17
rect -573 -34 -567 -32
rect -573 -36 -570 -34
rect -568 -36 -567 -34
rect -573 -41 -567 -36
rect -573 -43 -570 -41
rect -568 -43 -567 -41
rect -573 -45 -567 -43
rect -540 -24 -536 -19
rect -493 -13 -488 -11
rect -524 -24 -516 -23
rect -549 -25 -534 -24
rect -549 -27 -545 -25
rect -543 -27 -538 -25
rect -536 -27 -534 -25
rect -549 -28 -534 -27
rect -524 -26 -523 -24
rect -521 -25 -516 -24
rect -521 -26 -519 -25
rect -524 -27 -519 -26
rect -517 -27 -516 -25
rect -524 -29 -516 -27
rect -524 -32 -519 -29
rect -557 -36 -519 -32
rect -492 -35 -488 -13
rect -493 -37 -488 -35
rect -493 -39 -492 -37
rect -490 -39 -488 -37
rect -493 -44 -488 -39
rect -493 -46 -492 -44
rect -490 -46 -488 -44
rect -481 -16 -477 -7
rect -392 -9 -368 -8
rect -392 -11 -372 -9
rect -370 -11 -368 -9
rect -392 -12 -368 -11
rect -481 -18 -479 -16
rect -481 -34 -477 -18
rect -473 -16 -469 -15
rect -473 -18 -472 -16
rect -470 -18 -469 -16
rect -441 -16 -422 -15
rect -441 -17 -426 -16
rect -473 -23 -469 -18
rect -441 -19 -440 -17
rect -438 -18 -426 -17
rect -424 -18 -422 -16
rect -438 -19 -422 -18
rect -441 -20 -422 -19
rect -418 -17 -404 -16
rect -418 -19 -407 -17
rect -405 -19 -404 -17
rect -418 -20 -404 -19
rect -473 -25 -461 -23
rect -473 -27 -472 -25
rect -470 -27 -461 -25
rect -473 -29 -461 -27
rect -457 -25 -445 -23
rect -457 -27 -448 -25
rect -446 -27 -445 -25
rect -457 -29 -445 -27
rect -481 -36 -479 -34
rect -481 -39 -477 -36
rect -457 -37 -453 -29
rect -441 -32 -437 -20
rect -418 -24 -414 -20
rect -426 -25 -414 -24
rect -426 -27 -422 -25
rect -420 -27 -414 -25
rect -426 -28 -414 -27
rect -410 -25 -404 -24
rect -410 -27 -408 -25
rect -406 -27 -404 -25
rect -410 -32 -404 -27
rect -441 -34 -421 -32
rect -441 -36 -425 -34
rect -423 -36 -421 -34
rect -481 -41 -469 -39
rect -481 -43 -479 -41
rect -477 -43 -472 -41
rect -470 -43 -469 -41
rect -481 -45 -469 -43
rect -493 -48 -488 -46
rect -501 -49 -488 -48
rect -501 -51 -500 -49
rect -498 -51 -488 -49
rect -501 -52 -488 -51
rect -426 -41 -421 -36
rect -426 -43 -425 -41
rect -423 -43 -421 -41
rect -426 -45 -421 -43
rect -417 -37 -404 -32
rect -417 -42 -413 -37
rect -417 -44 -416 -42
rect -414 -44 -413 -42
rect -392 -40 -388 -12
rect -344 -19 -340 -17
rect -344 -21 -343 -19
rect -341 -21 -340 -19
rect -344 -22 -340 -21
rect -344 -24 -343 -22
rect -341 -24 -340 -22
rect -392 -41 -376 -40
rect -392 -43 -387 -41
rect -385 -43 -380 -41
rect -378 -43 -376 -41
rect -392 -44 -376 -43
rect -417 -45 -413 -44
rect -344 -38 -340 -24
rect -353 -39 -340 -38
rect -353 -41 -347 -39
rect -345 -41 -340 -39
rect -353 -44 -340 -41
rect -289 -23 -283 -16
rect -296 -24 -283 -23
rect -296 -26 -295 -24
rect -293 -26 -283 -24
rect -296 -29 -283 -26
rect -263 -16 -259 -7
rect -174 -9 -150 -8
rect -174 -11 -154 -9
rect -152 -11 -150 -9
rect -174 -12 -150 -11
rect -263 -18 -261 -16
rect -272 -24 -268 -23
rect -272 -26 -271 -24
rect -269 -26 -268 -24
rect -272 -30 -268 -26
rect -273 -32 -268 -30
rect -273 -34 -272 -32
rect -270 -34 -268 -32
rect -273 -36 -268 -34
rect -272 -40 -268 -36
rect -281 -41 -268 -40
rect -281 -43 -279 -41
rect -277 -43 -268 -41
rect -281 -45 -268 -43
rect -263 -34 -259 -18
rect -255 -16 -251 -15
rect -255 -18 -254 -16
rect -252 -18 -251 -16
rect -223 -16 -204 -15
rect -223 -17 -208 -16
rect -255 -23 -251 -18
rect -223 -19 -222 -17
rect -220 -18 -208 -17
rect -206 -18 -204 -16
rect -220 -19 -204 -18
rect -223 -20 -204 -19
rect -200 -17 -186 -16
rect -200 -19 -199 -17
rect -197 -19 -189 -17
rect -187 -19 -186 -17
rect -200 -20 -186 -19
rect -255 -25 -243 -23
rect -255 -27 -254 -25
rect -252 -27 -243 -25
rect -255 -29 -243 -27
rect -239 -25 -227 -23
rect -239 -27 -230 -25
rect -228 -27 -227 -25
rect -239 -29 -227 -27
rect -263 -36 -261 -34
rect -263 -39 -259 -36
rect -239 -37 -235 -29
rect -223 -32 -219 -20
rect -200 -24 -196 -20
rect -208 -25 -196 -24
rect -208 -27 -204 -25
rect -202 -27 -196 -25
rect -208 -28 -196 -27
rect -192 -25 -186 -24
rect -192 -27 -190 -25
rect -188 -27 -186 -25
rect -192 -32 -186 -27
rect -223 -34 -203 -32
rect -223 -36 -207 -34
rect -205 -36 -203 -34
rect -263 -41 -251 -39
rect -263 -43 -261 -41
rect -259 -43 -254 -41
rect -252 -43 -251 -41
rect -263 -45 -251 -43
rect -208 -41 -203 -36
rect -208 -43 -207 -41
rect -205 -43 -203 -41
rect -208 -45 -203 -43
rect -199 -37 -186 -32
rect -199 -42 -195 -37
rect -199 -44 -198 -42
rect -196 -44 -195 -42
rect -174 -40 -170 -12
rect -35 -9 -13 -8
rect -35 -11 -32 -9
rect -30 -11 -13 -9
rect -35 -12 -13 -11
rect 45 -9 50 -7
rect 45 -11 46 -9
rect 48 -11 50 -9
rect -126 -19 -122 -17
rect -126 -21 -125 -19
rect -123 -21 -122 -19
rect -126 -22 -122 -21
rect -126 -24 -125 -22
rect -123 -24 -122 -22
rect -174 -41 -158 -40
rect -174 -43 -166 -41
rect -164 -43 -162 -41
rect -160 -43 -158 -41
rect -174 -44 -158 -43
rect -199 -45 -195 -44
rect -126 -38 -122 -24
rect -135 -39 -122 -38
rect -135 -41 -129 -39
rect -127 -41 -122 -39
rect -135 -44 -122 -41
rect -71 -23 -65 -16
rect -78 -24 -65 -23
rect -78 -26 -77 -24
rect -75 -26 -65 -24
rect -78 -29 -65 -26
rect -54 -24 -50 -23
rect -54 -26 -53 -24
rect -51 -26 -50 -24
rect -54 -30 -50 -26
rect -55 -32 -50 -30
rect -55 -34 -54 -32
rect -52 -34 -50 -32
rect -55 -36 -50 -34
rect -54 -40 -50 -36
rect -63 -41 -50 -40
rect -63 -43 -61 -41
rect -59 -43 -50 -41
rect -63 -45 -50 -43
rect -35 -32 -31 -12
rect -2 -17 2 -15
rect -2 -19 -1 -17
rect 1 -19 2 -17
rect -35 -34 -29 -32
rect -35 -36 -32 -34
rect -30 -36 -29 -34
rect -35 -37 -29 -36
rect -35 -39 -33 -37
rect -31 -39 -29 -37
rect -35 -41 -29 -39
rect -35 -43 -32 -41
rect -30 -43 -29 -41
rect -35 -45 -29 -43
rect -2 -24 2 -19
rect 45 -13 50 -11
rect 14 -24 22 -23
rect -11 -25 4 -24
rect -11 -27 -7 -25
rect -5 -27 0 -25
rect 2 -27 4 -25
rect -11 -28 4 -27
rect 14 -26 15 -24
rect 17 -25 22 -24
rect 17 -26 19 -25
rect 14 -27 19 -26
rect 21 -27 22 -25
rect 14 -29 22 -27
rect 14 -32 19 -29
rect -19 -36 19 -32
rect 46 -35 50 -13
rect 45 -37 50 -35
rect 45 -39 46 -37
rect 48 -39 50 -37
rect 45 -44 50 -39
rect 45 -46 46 -44
rect 48 -46 50 -44
rect 45 -48 50 -46
rect 37 -52 50 -48
rect -584 -59 54 -58
rect -584 -61 -478 -59
rect -476 -61 -466 -59
rect -464 -61 -273 -59
rect -271 -61 -260 -59
rect -258 -61 -248 -59
rect -246 -61 -55 -59
rect -53 -61 54 -59
rect -584 -66 54 -61
rect -521 -71 13 -66
rect -521 -73 -514 -71
rect -512 -73 -502 -71
rect -500 -73 -309 -71
rect -307 -73 -294 -71
rect -292 -73 -282 -71
rect -280 -73 -89 -71
rect -87 -73 13 -71
rect -521 -74 13 -73
rect -517 -89 -505 -87
rect -517 -91 -515 -89
rect -513 -91 -505 -89
rect -517 -93 -505 -91
rect -462 -89 -457 -87
rect -462 -91 -461 -89
rect -459 -91 -457 -89
rect -517 -96 -513 -93
rect -517 -98 -515 -96
rect -517 -114 -513 -98
rect -493 -103 -489 -95
rect -462 -96 -457 -91
rect -477 -98 -461 -96
rect -459 -98 -457 -96
rect -477 -100 -457 -98
rect -453 -88 -449 -87
rect -453 -90 -452 -88
rect -450 -90 -449 -88
rect -453 -95 -449 -90
rect -428 -89 -412 -88
rect -428 -91 -416 -89
rect -414 -91 -412 -89
rect -428 -92 -412 -91
rect -453 -100 -440 -95
rect -509 -105 -497 -103
rect -509 -107 -508 -105
rect -506 -107 -497 -105
rect -509 -109 -497 -107
rect -493 -105 -481 -103
rect -493 -107 -484 -105
rect -482 -107 -481 -105
rect -493 -109 -481 -107
rect -517 -116 -515 -114
rect -517 -125 -513 -116
rect -509 -114 -505 -109
rect -509 -116 -508 -114
rect -506 -116 -505 -114
rect -477 -112 -473 -100
rect -462 -105 -450 -104
rect -462 -107 -458 -105
rect -456 -107 -450 -105
rect -462 -108 -450 -107
rect -446 -105 -440 -100
rect -446 -107 -444 -105
rect -442 -107 -440 -105
rect -446 -108 -440 -107
rect -454 -112 -450 -108
rect -477 -113 -458 -112
rect -477 -115 -476 -113
rect -474 -114 -458 -113
rect -474 -115 -462 -114
rect -509 -117 -505 -116
rect -477 -116 -462 -115
rect -460 -116 -458 -114
rect -454 -113 -440 -112
rect -454 -115 -443 -113
rect -441 -115 -440 -113
rect -454 -116 -440 -115
rect -477 -117 -458 -116
rect -428 -120 -424 -92
rect -389 -91 -376 -88
rect -389 -93 -383 -91
rect -381 -93 -376 -91
rect -389 -94 -376 -93
rect -428 -121 -404 -120
rect -428 -123 -408 -121
rect -406 -123 -404 -121
rect -428 -124 -404 -123
rect -380 -108 -376 -94
rect -380 -110 -379 -108
rect -377 -110 -376 -108
rect -380 -111 -376 -110
rect -380 -113 -379 -111
rect -377 -113 -376 -111
rect -380 -115 -376 -113
rect -317 -89 -304 -87
rect -317 -91 -315 -89
rect -313 -91 -304 -89
rect -317 -92 -304 -91
rect -308 -96 -304 -92
rect -332 -106 -319 -103
rect -332 -108 -331 -106
rect -329 -108 -319 -106
rect -332 -109 -319 -108
rect -325 -116 -319 -109
rect -309 -98 -304 -96
rect -309 -100 -308 -98
rect -306 -100 -304 -98
rect -309 -102 -304 -100
rect -308 -109 -304 -102
rect -297 -89 -285 -87
rect -297 -91 -295 -89
rect -293 -91 -285 -89
rect -297 -93 -285 -91
rect -4 -84 9 -80
rect -242 -89 -237 -87
rect -242 -91 -241 -89
rect -239 -91 -237 -89
rect -297 -96 -293 -93
rect -297 -98 -295 -96
rect -297 -114 -293 -98
rect -273 -103 -269 -95
rect -242 -96 -237 -91
rect -257 -98 -241 -96
rect -239 -98 -237 -96
rect -257 -100 -237 -98
rect -233 -88 -229 -87
rect -233 -90 -232 -88
rect -230 -90 -229 -88
rect -233 -95 -229 -90
rect -208 -89 -192 -88
rect -208 -91 -196 -89
rect -194 -91 -192 -89
rect -208 -92 -192 -91
rect -233 -100 -220 -95
rect -289 -105 -277 -103
rect -289 -107 -288 -105
rect -286 -107 -277 -105
rect -289 -109 -277 -107
rect -273 -105 -261 -103
rect -273 -107 -264 -105
rect -262 -107 -261 -105
rect -273 -109 -261 -107
rect -297 -116 -295 -114
rect -297 -125 -293 -116
rect -289 -114 -285 -109
rect -289 -116 -288 -114
rect -286 -116 -285 -114
rect -257 -112 -253 -100
rect -242 -105 -230 -104
rect -242 -107 -241 -105
rect -239 -107 -238 -105
rect -236 -107 -230 -105
rect -242 -108 -230 -107
rect -226 -105 -220 -100
rect -226 -107 -224 -105
rect -222 -107 -220 -105
rect -226 -108 -220 -107
rect -234 -112 -230 -108
rect -257 -113 -238 -112
rect -257 -115 -256 -113
rect -254 -114 -238 -113
rect -254 -115 -242 -114
rect -289 -117 -285 -116
rect -257 -116 -242 -115
rect -240 -116 -238 -114
rect -234 -113 -220 -112
rect -234 -115 -223 -113
rect -221 -115 -220 -113
rect -234 -116 -220 -115
rect -257 -117 -238 -116
rect -208 -120 -204 -92
rect -169 -91 -156 -88
rect -169 -93 -163 -91
rect -161 -93 -156 -91
rect -169 -94 -156 -93
rect -208 -121 -184 -120
rect -208 -123 -188 -121
rect -186 -123 -184 -121
rect -208 -124 -184 -123
rect -160 -108 -156 -94
rect -160 -110 -159 -108
rect -157 -110 -156 -108
rect -160 -111 -156 -110
rect -160 -113 -159 -111
rect -157 -113 -156 -111
rect -160 -115 -156 -113
rect -97 -89 -84 -87
rect -97 -91 -95 -89
rect -93 -91 -84 -89
rect -97 -92 -84 -91
rect -88 -96 -84 -92
rect -112 -106 -99 -103
rect -112 -108 -111 -106
rect -109 -108 -99 -106
rect -112 -109 -99 -108
rect -105 -116 -99 -109
rect -89 -98 -84 -96
rect -89 -100 -88 -98
rect -86 -100 -84 -98
rect -89 -102 -84 -100
rect -88 -109 -84 -102
rect -76 -89 -70 -87
rect 4 -86 9 -84
rect 4 -88 5 -86
rect 7 -88 9 -86
rect -76 -91 -73 -89
rect -71 -91 -70 -89
rect -76 -96 -70 -91
rect -76 -98 -73 -96
rect -71 -98 -70 -96
rect -76 -100 -70 -98
rect -76 -120 -72 -100
rect -60 -97 -22 -96
rect -60 -99 -34 -97
rect -32 -99 -22 -97
rect -60 -100 -22 -99
rect -27 -103 -22 -100
rect -52 -105 -37 -104
rect -52 -107 -51 -105
rect -49 -107 -48 -105
rect -46 -107 -41 -105
rect -39 -107 -37 -105
rect -52 -108 -37 -107
rect -27 -105 -19 -103
rect -27 -107 -22 -105
rect -20 -107 -19 -105
rect -43 -117 -39 -108
rect -27 -109 -19 -107
rect 4 -93 9 -88
rect 4 -95 5 -93
rect 7 -95 9 -93
rect 4 -97 9 -95
rect -76 -121 -54 -120
rect -76 -123 -73 -121
rect -71 -123 -54 -121
rect -76 -124 -54 -123
rect 5 -119 9 -97
rect 4 -121 9 -119
rect 4 -123 5 -121
rect 7 -123 9 -121
rect 4 -125 9 -123
rect -521 -131 13 -130
rect -521 -133 -514 -131
rect -512 -133 -502 -131
rect -500 -133 -480 -131
rect -478 -133 -426 -131
rect -424 -133 -364 -131
rect -362 -133 -309 -131
rect -307 -133 -294 -131
rect -292 -133 -282 -131
rect -280 -133 -260 -131
rect -258 -133 -206 -131
rect -204 -133 -144 -131
rect -142 -133 -89 -131
rect -87 -133 13 -131
rect -521 -138 13 -133
<< alu2 >>
rect -473 70 -469 71
rect -473 68 -472 70
rect -470 68 -469 70
rect -513 59 -509 60
rect -513 57 -512 59
rect -510 57 -509 59
rect -513 55 -509 57
rect -513 53 -512 55
rect -510 53 -509 55
rect -513 52 -509 53
rect -473 55 -469 68
rect -240 70 -236 71
rect -240 68 -239 70
rect -237 68 -236 70
rect -473 53 -472 55
rect -470 53 -469 55
rect -473 51 -469 53
rect -284 59 -280 60
rect -284 57 -283 59
rect -281 57 -280 59
rect -284 55 -280 57
rect -284 53 -283 55
rect -281 53 -280 55
rect -284 51 -280 53
rect -240 55 -236 68
rect -240 53 -239 55
rect -237 53 -236 55
rect -240 51 -236 53
rect -171 59 -167 60
rect -171 57 -170 59
rect -168 57 -167 59
rect -171 55 -167 57
rect -171 53 -170 55
rect -168 53 -167 55
rect -171 52 -167 53
rect -127 59 -123 61
rect -127 57 -126 59
rect -124 57 -123 59
rect -127 55 -123 57
rect -127 53 -126 55
rect -124 53 -123 55
rect -127 51 -123 53
rect -44 60 -40 61
rect -44 58 -43 60
rect -41 58 -40 60
rect -44 54 -40 58
rect -44 52 -43 54
rect -41 52 -40 54
rect -1 60 3 61
rect -1 58 0 60
rect 2 58 3 60
rect -1 55 3 58
rect -1 53 0 55
rect 2 53 3 55
rect -1 52 3 53
rect 82 60 86 61
rect 82 58 83 60
rect 85 58 86 60
rect 82 55 86 58
rect 82 53 83 55
rect 85 53 86 55
rect 82 52 86 53
rect -44 51 -40 52
rect -430 50 -426 51
rect -430 48 -429 50
rect -427 48 -426 50
rect -430 46 -426 48
rect -430 44 -429 46
rect -427 44 -426 46
rect -430 43 -426 44
rect -326 50 -322 51
rect -326 48 -325 50
rect -323 48 -322 50
rect -326 46 -322 48
rect -326 44 -325 46
rect -323 44 -322 46
rect -326 43 -322 44
rect -85 50 -81 51
rect -85 48 -84 50
rect -82 48 -81 50
rect -85 46 -81 48
rect -85 44 -84 46
rect -82 44 -81 46
rect -85 43 -81 44
rect 39 50 43 51
rect 39 48 40 50
rect 42 48 43 50
rect 39 46 43 48
rect 39 44 40 46
rect 42 44 43 46
rect 39 43 43 44
rect -521 37 -516 39
rect -521 35 -520 37
rect -518 35 -516 37
rect -540 21 -536 24
rect -540 19 -539 21
rect -537 19 -536 21
rect -540 -17 -536 19
rect -521 18 -516 35
rect -481 38 -476 39
rect -481 36 -480 38
rect -478 36 -476 38
rect -481 34 -476 36
rect -481 32 -479 34
rect -477 32 -476 34
rect -292 38 -287 39
rect -292 36 -291 38
rect -289 36 -287 38
rect -292 34 -287 36
rect -292 32 -290 34
rect -288 32 -287 34
rect -481 31 -476 32
rect -438 29 -433 31
rect -438 27 -436 29
rect -434 27 -433 29
rect -521 16 -520 18
rect -518 16 -516 18
rect -521 15 -516 16
rect -505 21 -500 24
rect -505 19 -503 21
rect -501 19 -500 21
rect -540 -19 -539 -17
rect -537 -19 -536 -17
rect -540 -21 -536 -19
rect -524 -10 -519 -9
rect -524 -12 -522 -10
rect -520 -12 -519 -10
rect -524 -24 -519 -12
rect -505 -10 -500 19
rect -461 21 -457 24
rect -461 19 -460 21
rect -458 19 -457 21
rect -505 -12 -503 -10
rect -501 -12 -500 -10
rect -505 -13 -500 -12
rect -473 -11 -469 -10
rect -473 -13 -472 -11
rect -470 -13 -469 -11
rect -473 -16 -469 -13
rect -473 -18 -472 -16
rect -470 -18 -469 -16
rect -473 -19 -469 -18
rect -524 -26 -523 -24
rect -521 -26 -519 -24
rect -524 -28 -519 -26
rect -473 -41 -469 -39
rect -473 -43 -472 -41
rect -470 -43 -469 -41
rect -501 -49 -497 -48
rect -501 -51 -500 -49
rect -498 -51 -497 -49
rect -501 -97 -497 -51
rect -473 -82 -469 -43
rect -461 -59 -457 19
rect -438 7 -433 27
rect -334 30 -329 32
rect -292 31 -287 32
rect -93 38 -88 39
rect -93 36 -92 38
rect -90 36 -88 38
rect -93 34 -88 36
rect -93 32 -92 34
rect -90 32 -88 34
rect -93 31 -88 32
rect -9 38 -4 39
rect -9 36 -8 38
rect -6 36 -4 38
rect -9 34 -4 36
rect -9 32 -8 34
rect -6 32 -4 34
rect -9 31 -4 32
rect -334 28 -333 30
rect -331 28 -329 30
rect -438 5 -437 7
rect -435 5 -433 7
rect -438 4 -433 5
rect -354 21 -350 24
rect -354 19 -353 21
rect -351 19 -350 21
rect -441 -11 -437 -10
rect -441 -13 -440 -11
rect -438 -13 -437 -11
rect -441 -17 -437 -13
rect -441 -19 -440 -17
rect -438 -19 -437 -17
rect -441 -20 -437 -19
rect -408 -13 -404 -12
rect -408 -15 -407 -13
rect -405 -15 -404 -13
rect -408 -17 -404 -15
rect -354 -13 -350 19
rect -334 18 -329 28
rect -272 30 -268 31
rect -272 28 -271 30
rect -269 28 -268 30
rect -334 16 -332 18
rect -330 16 -329 18
rect -334 15 -329 16
rect -316 21 -312 24
rect -316 19 -315 21
rect -313 19 -312 21
rect -354 -15 -353 -13
rect -351 -15 -350 -13
rect -354 -16 -350 -15
rect -344 -15 -340 -13
rect -408 -19 -407 -17
rect -405 -19 -404 -17
rect -408 -20 -404 -19
rect -344 -17 -343 -15
rect -341 -17 -340 -15
rect -344 -22 -340 -17
rect -450 -25 -445 -23
rect -344 -24 -343 -22
rect -341 -24 -340 -22
rect -344 -25 -340 -24
rect -450 -27 -448 -25
rect -446 -27 -445 -25
rect -450 -33 -445 -27
rect -450 -35 -448 -33
rect -446 -35 -445 -33
rect -450 -36 -445 -35
rect -316 -33 -312 19
rect -316 -35 -315 -33
rect -313 -35 -312 -33
rect -316 -36 -312 -35
rect -296 -24 -290 -23
rect -296 -26 -295 -24
rect -293 -26 -290 -24
rect -296 -33 -290 -26
rect -272 -24 -268 28
rect -248 30 -243 31
rect -248 28 -247 30
rect -245 28 -243 30
rect -248 26 -243 28
rect -248 24 -247 26
rect -245 24 -243 26
rect -179 30 -174 31
rect -179 28 -178 30
rect -176 28 -174 30
rect -179 26 -174 28
rect -179 24 -178 26
rect -176 24 -174 26
rect -248 23 -243 24
rect -200 21 -196 24
rect -179 23 -174 24
rect -135 30 -130 31
rect -135 28 -134 30
rect -132 28 -130 30
rect -200 19 -199 21
rect -197 19 -196 21
rect -255 -11 -251 -10
rect -255 -13 -254 -11
rect -252 -13 -251 -11
rect -255 -16 -251 -13
rect -255 -18 -254 -16
rect -252 -18 -251 -16
rect -255 -19 -251 -18
rect -223 -11 -219 -10
rect -223 -13 -222 -11
rect -220 -13 -219 -11
rect -223 -17 -219 -13
rect -223 -19 -222 -17
rect -220 -19 -219 -17
rect -223 -20 -219 -19
rect -200 -17 -196 19
rect -151 22 -147 23
rect -151 20 -150 22
rect -148 20 -147 22
rect -200 -19 -199 -17
rect -197 -19 -196 -17
rect -200 -21 -196 -19
rect -190 -13 -186 -12
rect -190 -15 -189 -13
rect -187 -15 -186 -13
rect -190 -17 -186 -15
rect -190 -19 -189 -17
rect -187 -19 -186 -17
rect -190 -20 -186 -19
rect -272 -26 -271 -24
rect -269 -26 -268 -24
rect -272 -27 -268 -26
rect -232 -25 -227 -23
rect -232 -27 -230 -25
rect -228 -27 -227 -25
rect -296 -35 -294 -33
rect -292 -35 -290 -33
rect -296 -36 -290 -35
rect -232 -33 -227 -27
rect -232 -35 -230 -33
rect -228 -35 -227 -33
rect -232 -36 -227 -35
rect -388 -41 -384 -40
rect -417 -42 -413 -41
rect -417 -44 -416 -42
rect -414 -44 -413 -42
rect -417 -48 -413 -44
rect -417 -50 -416 -48
rect -414 -50 -413 -48
rect -417 -51 -413 -50
rect -388 -43 -387 -41
rect -385 -43 -384 -41
rect -461 -61 -460 -59
rect -458 -61 -457 -59
rect -461 -62 -457 -61
rect -444 -59 -440 -54
rect -444 -61 -443 -59
rect -441 -61 -440 -59
rect -473 -84 -472 -82
rect -470 -84 -469 -82
rect -473 -85 -469 -84
rect -453 -82 -449 -81
rect -453 -84 -452 -82
rect -450 -84 -449 -82
rect -453 -88 -449 -84
rect -453 -90 -452 -88
rect -450 -90 -449 -88
rect -453 -91 -449 -90
rect -501 -99 -500 -97
rect -498 -99 -497 -97
rect -501 -100 -497 -99
rect -486 -97 -481 -96
rect -486 -99 -484 -97
rect -482 -99 -481 -97
rect -486 -105 -481 -99
rect -486 -107 -484 -105
rect -482 -107 -481 -105
rect -486 -109 -481 -107
rect -477 -113 -473 -112
rect -509 -114 -505 -113
rect -509 -116 -508 -114
rect -506 -116 -505 -114
rect -509 -119 -505 -116
rect -509 -121 -508 -119
rect -506 -121 -505 -119
rect -509 -122 -505 -121
rect -477 -115 -476 -113
rect -474 -115 -473 -113
rect -477 -119 -473 -115
rect -477 -121 -476 -119
rect -474 -121 -473 -119
rect -444 -113 -440 -61
rect -388 -61 -384 -43
rect -280 -41 -276 -40
rect -280 -43 -279 -41
rect -277 -43 -276 -41
rect -280 -48 -276 -43
rect -280 -50 -279 -48
rect -277 -50 -276 -48
rect -280 -51 -276 -50
rect -255 -41 -251 -39
rect -167 -41 -163 -40
rect -255 -43 -254 -41
rect -252 -43 -251 -41
rect -388 -63 -387 -61
rect -385 -63 -384 -61
rect -388 -64 -384 -63
rect -266 -61 -261 -60
rect -266 -63 -264 -61
rect -262 -63 -261 -61
rect -316 -82 -312 -81
rect -316 -84 -315 -82
rect -313 -84 -312 -82
rect -316 -89 -312 -84
rect -316 -91 -315 -89
rect -313 -91 -312 -89
rect -316 -92 -312 -91
rect -332 -97 -326 -96
rect -332 -99 -330 -97
rect -328 -99 -326 -97
rect -332 -106 -326 -99
rect -444 -115 -443 -113
rect -441 -115 -440 -113
rect -444 -117 -440 -115
rect -444 -119 -443 -117
rect -441 -119 -440 -117
rect -380 -108 -376 -107
rect -380 -110 -379 -108
rect -377 -110 -376 -108
rect -332 -108 -331 -106
rect -329 -108 -326 -106
rect -332 -109 -326 -108
rect -266 -97 -261 -63
rect -255 -82 -251 -43
rect -199 -42 -195 -41
rect -199 -44 -198 -42
rect -196 -44 -195 -42
rect -199 -48 -195 -44
rect -199 -50 -198 -48
rect -196 -50 -195 -48
rect -199 -51 -195 -50
rect -167 -43 -166 -41
rect -164 -43 -163 -41
rect -167 -59 -163 -43
rect -167 -61 -166 -59
rect -164 -61 -163 -59
rect -167 -62 -163 -61
rect -255 -84 -254 -82
rect -252 -84 -251 -82
rect -255 -85 -251 -84
rect -242 -82 -238 -81
rect -242 -84 -241 -82
rect -239 -84 -238 -82
rect -266 -99 -264 -97
rect -262 -99 -261 -97
rect -266 -105 -261 -99
rect -266 -107 -264 -105
rect -262 -107 -261 -105
rect -266 -109 -261 -107
rect -242 -105 -238 -84
rect -233 -82 -229 -81
rect -233 -84 -232 -82
rect -230 -84 -229 -82
rect -233 -88 -229 -84
rect -151 -82 -147 20
rect -135 8 -130 28
rect -52 30 -47 31
rect -52 28 -51 30
rect -49 28 -47 30
rect -135 6 -134 8
rect -132 6 -130 8
rect -135 4 -130 6
rect -117 21 -113 22
rect -117 19 -116 21
rect -114 19 -113 21
rect -126 -15 -122 -13
rect -126 -17 -125 -15
rect -123 -17 -122 -15
rect -126 -22 -122 -17
rect -126 -24 -125 -22
rect -123 -24 -122 -22
rect -126 -25 -122 -24
rect -117 -33 -113 19
rect -69 21 -64 23
rect -69 19 -68 21
rect -66 19 -64 21
rect -69 -9 -64 19
rect -52 18 -47 28
rect 32 29 36 31
rect 32 27 33 29
rect 35 27 36 29
rect 32 26 36 27
rect 32 24 33 26
rect 35 24 36 26
rect -52 16 -50 18
rect -48 16 -47 18
rect -52 15 -47 16
rect -26 21 -21 24
rect 32 23 36 24
rect 75 29 79 31
rect 75 27 76 29
rect 78 27 79 29
rect 75 26 79 27
rect 75 24 76 26
rect 78 24 79 26
rect 75 23 79 24
rect -26 19 -25 21
rect -23 19 -21 21
rect -69 -11 -68 -9
rect -66 -11 -64 -9
rect -69 -12 -64 -11
rect -54 -9 -50 -8
rect -54 -11 -53 -9
rect -51 -11 -50 -9
rect -117 -35 -116 -33
rect -114 -35 -113 -33
rect -117 -36 -113 -35
rect -78 -24 -72 -23
rect -78 -26 -77 -24
rect -75 -26 -72 -24
rect -78 -33 -72 -26
rect -54 -24 -50 -11
rect -26 -9 -21 19
rect 14 21 19 22
rect 14 19 15 21
rect 17 19 19 21
rect -26 -11 -25 -9
rect -23 -11 -21 -9
rect -26 -12 -21 -11
rect -2 -9 2 -8
rect -2 -11 -1 -9
rect 1 -11 2 -9
rect -2 -17 2 -11
rect -2 -19 -1 -17
rect 1 -19 2 -17
rect -2 -20 2 -19
rect -54 -26 -53 -24
rect -51 -26 -50 -24
rect -54 -27 -50 -26
rect 14 -24 19 19
rect 14 -26 15 -24
rect 17 -26 19 -24
rect 14 -27 19 -26
rect -78 -35 -76 -33
rect -74 -35 -72 -33
rect -78 -36 -72 -35
rect -35 -37 -29 -32
rect -35 -39 -33 -37
rect -31 -39 -29 -37
rect -62 -41 -58 -40
rect -62 -43 -61 -41
rect -59 -43 -58 -41
rect -62 -48 -58 -43
rect -62 -50 -61 -48
rect -59 -50 -58 -48
rect -62 -51 -58 -50
rect -52 -59 -48 -58
rect -52 -61 -51 -59
rect -49 -61 -48 -59
rect -151 -84 -150 -82
rect -148 -84 -147 -82
rect -151 -85 -147 -84
rect -96 -82 -92 -81
rect -96 -84 -95 -82
rect -93 -84 -92 -82
rect -233 -90 -232 -88
rect -230 -90 -229 -88
rect -233 -91 -229 -90
rect -96 -89 -92 -84
rect -96 -91 -95 -89
rect -93 -91 -92 -89
rect -96 -92 -92 -91
rect -242 -107 -241 -105
rect -239 -107 -238 -105
rect -112 -97 -106 -96
rect -112 -99 -110 -97
rect -108 -99 -106 -97
rect -112 -106 -106 -99
rect -242 -108 -238 -107
rect -160 -108 -156 -107
rect -380 -115 -376 -110
rect -160 -110 -159 -108
rect -157 -110 -156 -108
rect -112 -108 -111 -106
rect -109 -108 -106 -106
rect -52 -105 -48 -61
rect -35 -97 -29 -39
rect -35 -99 -34 -97
rect -32 -99 -29 -97
rect -35 -100 -29 -99
rect -52 -107 -51 -105
rect -49 -107 -48 -105
rect -52 -108 -48 -107
rect -112 -109 -106 -108
rect -257 -113 -253 -112
rect -380 -117 -379 -115
rect -377 -117 -376 -115
rect -380 -119 -376 -117
rect -289 -114 -285 -113
rect -289 -116 -288 -114
rect -286 -116 -285 -114
rect -289 -119 -285 -116
rect -444 -120 -440 -119
rect -477 -122 -473 -121
rect -289 -121 -288 -119
rect -286 -121 -285 -119
rect -289 -122 -285 -121
rect -257 -115 -256 -113
rect -254 -115 -253 -113
rect -257 -119 -253 -115
rect -257 -121 -256 -119
rect -254 -121 -253 -119
rect -224 -113 -220 -112
rect -224 -115 -223 -113
rect -221 -115 -220 -113
rect -224 -117 -220 -115
rect -224 -119 -223 -117
rect -221 -119 -220 -117
rect -160 -115 -156 -110
rect -160 -117 -159 -115
rect -157 -117 -156 -115
rect -160 -119 -156 -117
rect -224 -120 -220 -119
rect -257 -122 -253 -121
<< alu3 >>
rect -473 70 -236 71
rect -473 68 -472 70
rect -470 68 -239 70
rect -237 68 -236 70
rect -473 67 -236 68
rect -127 60 86 61
rect -513 59 -167 60
rect -513 57 -512 59
rect -510 57 -283 59
rect -281 57 -170 59
rect -168 57 -167 59
rect -513 56 -167 57
rect -127 59 -43 60
rect -127 57 -126 59
rect -124 58 -43 59
rect -41 58 0 60
rect 2 58 83 60
rect 85 58 86 60
rect -124 57 86 58
rect -127 56 86 57
rect -430 46 43 47
rect -430 44 -429 46
rect -427 44 -325 46
rect -323 44 -84 46
rect -82 44 40 46
rect 42 44 43 46
rect -430 43 43 44
rect -481 34 -4 35
rect -481 32 -479 34
rect -477 32 -290 34
rect -288 32 -92 34
rect -90 32 -8 34
rect -6 32 -4 34
rect -481 31 -4 32
rect -248 26 79 27
rect -248 24 -247 26
rect -245 24 -178 26
rect -176 24 33 26
rect 35 24 76 26
rect 78 24 79 26
rect -248 23 79 24
rect -521 18 -47 19
rect -521 16 -520 18
rect -518 16 -332 18
rect -330 16 -50 18
rect -48 16 -47 18
rect -521 15 -47 16
rect -438 8 -130 9
rect -438 7 -134 8
rect -438 5 -437 7
rect -435 6 -134 7
rect -132 6 -130 8
rect -435 5 -130 6
rect -438 4 -130 5
rect -69 -9 -50 -8
rect -524 -10 -500 -9
rect -524 -12 -522 -10
rect -520 -12 -503 -10
rect -501 -12 -500 -10
rect -524 -13 -500 -12
rect -473 -11 -436 -10
rect -473 -13 -472 -11
rect -470 -13 -440 -11
rect -438 -13 -436 -11
rect -255 -11 -218 -10
rect -473 -14 -436 -13
rect -408 -13 -340 -12
rect -408 -15 -407 -13
rect -405 -15 -353 -13
rect -351 -15 -340 -13
rect -255 -13 -254 -11
rect -252 -13 -222 -11
rect -220 -13 -218 -11
rect -69 -11 -68 -9
rect -66 -11 -53 -9
rect -51 -11 -50 -9
rect -69 -12 -50 -11
rect -26 -9 2 -8
rect -26 -11 -25 -9
rect -23 -11 -1 -9
rect 1 -11 2 -9
rect -26 -12 2 -11
rect -255 -14 -218 -13
rect -190 -13 -122 -12
rect -408 -16 -343 -15
rect -344 -17 -343 -16
rect -341 -17 -340 -15
rect -190 -15 -189 -13
rect -187 -15 -122 -13
rect -190 -16 -125 -15
rect -344 -18 -340 -17
rect -126 -17 -125 -16
rect -123 -17 -122 -15
rect -126 -18 -122 -17
rect -450 -33 -290 -32
rect -450 -35 -448 -33
rect -446 -35 -315 -33
rect -313 -35 -294 -33
rect -292 -35 -290 -33
rect -450 -36 -290 -35
rect -232 -33 -72 -32
rect -232 -35 -230 -33
rect -228 -35 -116 -33
rect -114 -35 -76 -33
rect -74 -35 -72 -33
rect -232 -36 -72 -35
rect -417 -48 -276 -47
rect -417 -50 -416 -48
rect -414 -50 -279 -48
rect -277 -50 -276 -48
rect -417 -51 -276 -50
rect -199 -48 -58 -47
rect -199 -50 -198 -48
rect -196 -50 -61 -48
rect -59 -50 -58 -48
rect -199 -51 -58 -50
rect -461 -59 -440 -58
rect -461 -61 -460 -59
rect -458 -61 -443 -59
rect -441 -61 -440 -59
rect -167 -59 -48 -58
rect -461 -62 -440 -61
rect -388 -61 -261 -60
rect -388 -63 -387 -61
rect -385 -63 -264 -61
rect -262 -63 -261 -61
rect -167 -61 -166 -59
rect -164 -61 -51 -59
rect -49 -61 -48 -59
rect -167 -62 -48 -61
rect -388 -64 -261 -63
rect -473 -82 -312 -81
rect -473 -84 -472 -82
rect -470 -84 -452 -82
rect -450 -84 -315 -82
rect -313 -84 -312 -82
rect -473 -85 -312 -84
rect -255 -82 -238 -81
rect -255 -84 -254 -82
rect -252 -84 -241 -82
rect -239 -84 -238 -82
rect -255 -85 -238 -84
rect -233 -82 -92 -81
rect -233 -84 -232 -82
rect -230 -84 -150 -82
rect -148 -84 -95 -82
rect -93 -84 -92 -82
rect -233 -85 -92 -84
rect -501 -97 -326 -96
rect -501 -99 -500 -97
rect -498 -99 -484 -97
rect -482 -99 -330 -97
rect -328 -99 -326 -97
rect -501 -100 -326 -99
rect -266 -97 -106 -96
rect -266 -99 -264 -97
rect -262 -99 -110 -97
rect -108 -99 -106 -97
rect -266 -100 -106 -99
rect -380 -115 -376 -114
rect -380 -116 -379 -115
rect -444 -117 -379 -116
rect -377 -117 -376 -115
rect -160 -115 -156 -114
rect -160 -116 -159 -115
rect -509 -119 -472 -118
rect -509 -121 -508 -119
rect -506 -121 -476 -119
rect -474 -121 -472 -119
rect -444 -119 -443 -117
rect -441 -119 -376 -117
rect -224 -117 -159 -116
rect -157 -117 -156 -115
rect -444 -120 -376 -119
rect -289 -119 -252 -118
rect -509 -122 -472 -121
rect -289 -121 -288 -119
rect -286 -121 -256 -119
rect -254 -121 -252 -119
rect -224 -119 -223 -117
rect -221 -119 -156 -117
rect -224 -120 -156 -119
rect -289 -122 -252 -121
<< ptie >>
rect -544 12 -538 14
rect -544 10 -542 12
rect -540 10 -538 12
rect -544 8 -538 10
rect -504 12 -498 14
rect -504 10 -502 12
rect -500 10 -498 12
rect -504 8 -498 10
rect -461 12 -455 14
rect -461 10 -459 12
rect -457 10 -455 12
rect -461 8 -455 10
rect -357 12 -351 14
rect -357 10 -355 12
rect -353 10 -351 12
rect -357 8 -351 10
rect -315 12 -309 14
rect -315 10 -313 12
rect -311 10 -309 12
rect -315 8 -309 10
rect -271 12 -265 14
rect -271 10 -269 12
rect -267 10 -265 12
rect -271 8 -265 10
rect -202 12 -196 14
rect -202 10 -200 12
rect -198 10 -196 12
rect -202 8 -196 10
rect -158 12 -152 14
rect -158 10 -156 12
rect -154 10 -152 12
rect -158 8 -152 10
rect -116 12 -110 14
rect -116 10 -114 12
rect -112 10 -110 12
rect -116 8 -110 10
rect -75 12 -69 14
rect -75 10 -73 12
rect -71 10 -69 12
rect -75 8 -69 10
rect -32 12 -26 14
rect -32 10 -30 12
rect -28 10 -26 12
rect -32 8 -26 10
rect 8 12 14 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 51 12 57 14
rect 51 10 53 12
rect 55 10 57 12
rect 51 8 57 10
rect -480 1 -462 3
rect -480 -1 -478 1
rect -476 -1 -466 1
rect -464 -1 -462 1
rect -480 -3 -462 -1
rect -275 1 -269 3
rect -275 -1 -273 1
rect -271 -1 -269 1
rect -275 -3 -269 -1
rect -262 1 -244 3
rect -262 -1 -260 1
rect -258 -1 -248 1
rect -246 -1 -244 1
rect -262 -3 -244 -1
rect -57 1 -51 3
rect -57 -1 -55 1
rect -53 -1 -51 1
rect -57 -3 -51 -1
rect -516 -131 -498 -129
rect -516 -133 -514 -131
rect -512 -133 -502 -131
rect -500 -133 -498 -131
rect -516 -135 -498 -133
rect -311 -131 -305 -129
rect -311 -133 -309 -131
rect -307 -133 -305 -131
rect -311 -135 -305 -133
rect -296 -131 -278 -129
rect -296 -133 -294 -131
rect -292 -133 -282 -131
rect -280 -133 -278 -131
rect -296 -135 -278 -133
rect -91 -131 -85 -129
rect -91 -133 -89 -131
rect -87 -133 -85 -131
rect -91 -135 -85 -133
<< ntie >>
rect -544 72 -538 74
rect -544 70 -542 72
rect -540 70 -538 72
rect -544 68 -538 70
rect -504 72 -498 74
rect -504 70 -502 72
rect -500 70 -498 72
rect -504 68 -498 70
rect -461 72 -455 74
rect -461 70 -459 72
rect -457 70 -455 72
rect -461 68 -455 70
rect -357 72 -351 74
rect -357 70 -355 72
rect -353 70 -351 72
rect -357 68 -351 70
rect -315 72 -309 74
rect -315 70 -313 72
rect -311 70 -309 72
rect -315 68 -309 70
rect -271 72 -265 74
rect -271 70 -269 72
rect -267 70 -265 72
rect -271 68 -265 70
rect -202 72 -196 74
rect -202 70 -200 72
rect -198 70 -196 72
rect -202 68 -196 70
rect -158 72 -152 74
rect -158 70 -156 72
rect -154 70 -152 72
rect -158 68 -152 70
rect -116 72 -110 74
rect -116 70 -114 72
rect -112 70 -110 72
rect -116 68 -110 70
rect -75 72 -69 74
rect -75 70 -73 72
rect -71 70 -69 72
rect -75 68 -69 70
rect -32 72 -26 74
rect -32 70 -30 72
rect -28 70 -26 72
rect -32 68 -26 70
rect 8 72 14 74
rect 8 70 10 72
rect 12 70 14 72
rect 8 68 14 70
rect 51 72 57 74
rect 51 70 53 72
rect 55 70 57 72
rect 51 68 57 70
rect -480 -59 -462 -57
rect -480 -61 -478 -59
rect -476 -61 -466 -59
rect -464 -61 -462 -59
rect -480 -63 -462 -61
rect -275 -59 -269 -57
rect -275 -61 -273 -59
rect -271 -61 -269 -59
rect -275 -63 -269 -61
rect -262 -59 -244 -57
rect -262 -61 -260 -59
rect -258 -61 -248 -59
rect -246 -61 -244 -59
rect -262 -63 -244 -61
rect -57 -59 -51 -57
rect -57 -61 -55 -59
rect -53 -61 -51 -59
rect -57 -63 -51 -61
rect -516 -71 -498 -69
rect -516 -73 -514 -71
rect -512 -73 -502 -71
rect -500 -73 -498 -71
rect -311 -71 -305 -69
rect -516 -75 -498 -73
rect -311 -73 -309 -71
rect -307 -73 -305 -71
rect -311 -75 -305 -73
rect -296 -71 -278 -69
rect -296 -73 -294 -71
rect -292 -73 -282 -71
rect -280 -73 -278 -71
rect -91 -71 -85 -69
rect -296 -75 -278 -73
rect -91 -73 -89 -71
rect -87 -73 -85 -71
rect -91 -75 -85 -73
<< nmos >>
rect -538 20 -536 29
rect -525 18 -523 29
rect -518 18 -516 29
rect -498 20 -496 29
rect -485 18 -483 29
rect -478 18 -476 29
rect -455 20 -453 29
rect -442 18 -440 29
rect -435 18 -433 29
rect -351 20 -349 29
rect -338 18 -336 29
rect -331 18 -329 29
rect -309 20 -307 29
rect -296 18 -294 29
rect -289 18 -287 29
rect -265 20 -263 29
rect -252 18 -250 29
rect -245 18 -243 29
rect -196 20 -194 29
rect -183 18 -181 29
rect -176 18 -174 29
rect -152 20 -150 29
rect -139 18 -137 29
rect -132 18 -130 29
rect -110 20 -108 29
rect -97 18 -95 29
rect -90 18 -88 29
rect -69 20 -67 29
rect -56 18 -54 29
rect -49 18 -47 29
rect -26 20 -24 29
rect -13 18 -11 29
rect -6 18 -4 29
rect 14 20 16 29
rect 27 18 29 29
rect 34 18 36 29
rect 57 20 59 29
rect 70 18 72 29
rect 77 18 79 29
rect -565 -14 -563 0
rect -554 -20 -552 0
rect -547 -20 -545 0
rect -527 -20 -525 -6
rect -517 -20 -515 -6
rect -507 -13 -505 -3
rect -497 -13 -495 0
rect -474 -20 -472 -11
rect -450 -18 -448 -6
rect -438 -20 -436 -8
rect -431 -20 -429 -8
rect -421 -20 -419 -8
rect -411 -20 -409 -8
rect -384 -14 -382 -1
rect -377 -14 -375 -1
rect -367 -14 -365 -1
rect -357 -19 -355 -6
rect -345 -14 -343 -3
rect -322 -14 -320 -1
rect -315 -14 -313 -1
rect -305 -14 -303 -1
rect -295 -19 -293 -6
rect -284 -20 -282 -9
rect -256 -20 -254 -11
rect -232 -18 -230 -6
rect -220 -20 -218 -8
rect -213 -20 -211 -8
rect -203 -20 -201 -8
rect -193 -20 -191 -8
rect -166 -14 -164 -1
rect -159 -14 -157 -1
rect -149 -14 -147 -1
rect -139 -19 -137 -6
rect -127 -14 -125 -3
rect -104 -14 -102 -1
rect -97 -14 -95 -1
rect -87 -14 -85 -1
rect -77 -19 -75 -6
rect -66 -20 -64 -9
rect -27 -14 -25 0
rect -16 -20 -14 0
rect -9 -20 -7 0
rect 11 -20 13 -6
rect 21 -20 23 -6
rect 31 -13 33 -3
rect 41 -13 43 0
rect -510 -121 -508 -112
rect -486 -126 -484 -114
rect -474 -124 -472 -112
rect -467 -124 -465 -112
rect -457 -124 -455 -112
rect -447 -124 -445 -112
rect -420 -131 -418 -118
rect -413 -131 -411 -118
rect -403 -131 -401 -118
rect -393 -126 -391 -113
rect -381 -129 -379 -118
rect -358 -131 -356 -118
rect -351 -131 -349 -118
rect -341 -131 -339 -118
rect -331 -126 -329 -113
rect -320 -123 -318 -112
rect -290 -121 -288 -112
rect -266 -126 -264 -114
rect -254 -124 -252 -112
rect -247 -124 -245 -112
rect -237 -124 -235 -112
rect -227 -124 -225 -112
rect -200 -131 -198 -118
rect -193 -131 -191 -118
rect -183 -131 -181 -118
rect -173 -126 -171 -113
rect -161 -129 -159 -118
rect -138 -131 -136 -118
rect -131 -131 -129 -118
rect -121 -131 -119 -118
rect -111 -126 -109 -113
rect -100 -123 -98 -112
rect -68 -132 -66 -118
rect -57 -132 -55 -112
rect -50 -132 -48 -112
rect -30 -126 -28 -112
rect -20 -126 -18 -112
rect -10 -129 -8 -119
rect 0 -132 2 -119
<< pmos >>
rect -538 44 -536 62
rect -528 51 -526 64
rect -518 51 -516 64
rect -498 44 -496 62
rect -488 51 -486 64
rect -478 51 -476 64
rect -455 44 -453 62
rect -445 51 -443 64
rect -435 51 -433 64
rect -351 44 -349 62
rect -341 51 -339 64
rect -331 51 -329 64
rect -309 44 -307 62
rect -299 51 -297 64
rect -289 51 -287 64
rect -265 44 -263 62
rect -255 51 -253 64
rect -245 51 -243 64
rect -196 44 -194 62
rect -186 51 -184 64
rect -176 51 -174 64
rect -152 44 -150 62
rect -142 51 -140 64
rect -132 51 -130 64
rect -110 44 -108 62
rect -100 51 -98 64
rect -90 51 -88 64
rect -69 44 -67 62
rect -59 51 -57 64
rect -49 51 -47 64
rect -26 44 -24 62
rect -16 51 -14 64
rect -6 51 -4 64
rect 14 44 16 62
rect 24 51 26 64
rect 34 51 36 64
rect 57 44 59 62
rect 67 51 69 64
rect 77 51 79 64
rect -565 -60 -563 -32
rect -555 -60 -553 -32
rect -545 -60 -543 -32
rect -527 -57 -525 -32
rect -520 -57 -518 -32
rect -510 -48 -508 -35
rect -497 -60 -495 -35
rect -474 -50 -472 -32
rect -447 -59 -445 -32
rect -437 -59 -435 -32
rect -430 -59 -428 -32
rect -420 -59 -418 -32
rect -410 -59 -408 -32
rect -385 -60 -383 -32
rect -375 -60 -373 -32
rect -365 -60 -363 -32
rect -355 -60 -353 -46
rect -345 -60 -343 -46
rect -325 -60 -323 -32
rect -315 -60 -313 -32
rect -305 -60 -303 -32
rect -294 -53 -292 -39
rect -284 -53 -282 -39
rect -256 -50 -254 -32
rect -229 -59 -227 -32
rect -219 -59 -217 -32
rect -212 -59 -210 -32
rect -202 -59 -200 -32
rect -192 -59 -190 -32
rect -167 -60 -165 -32
rect -157 -60 -155 -32
rect -147 -60 -145 -32
rect -137 -60 -135 -46
rect -127 -60 -125 -46
rect -107 -60 -105 -32
rect -97 -60 -95 -32
rect -87 -60 -85 -32
rect -76 -53 -74 -39
rect -66 -53 -64 -39
rect -27 -60 -25 -32
rect -17 -60 -15 -32
rect -7 -60 -5 -32
rect 11 -57 13 -32
rect 18 -57 20 -32
rect 28 -48 30 -35
rect 41 -60 43 -35
rect -510 -100 -508 -82
rect -483 -100 -481 -73
rect -473 -100 -471 -73
rect -466 -100 -464 -73
rect -456 -100 -454 -73
rect -446 -100 -444 -73
rect -421 -100 -419 -72
rect -411 -100 -409 -72
rect -401 -100 -399 -72
rect -391 -86 -389 -72
rect -381 -86 -379 -72
rect -361 -100 -359 -72
rect -351 -100 -349 -72
rect -341 -100 -339 -72
rect -330 -93 -328 -79
rect -320 -93 -318 -79
rect -290 -100 -288 -82
rect -263 -100 -261 -73
rect -253 -100 -251 -73
rect -246 -100 -244 -73
rect -236 -100 -234 -73
rect -226 -100 -224 -73
rect -201 -100 -199 -72
rect -191 -100 -189 -72
rect -181 -100 -179 -72
rect -171 -86 -169 -72
rect -161 -86 -159 -72
rect -141 -100 -139 -72
rect -131 -100 -129 -72
rect -121 -100 -119 -72
rect -110 -93 -108 -79
rect -100 -93 -98 -79
rect -68 -100 -66 -72
rect -58 -100 -56 -72
rect -48 -100 -46 -72
rect -30 -100 -28 -75
rect -23 -100 -21 -75
rect -13 -97 -11 -84
rect 0 -97 2 -72
<< polyct0 >>
rect -536 36 -534 38
rect -496 36 -494 38
rect -453 36 -451 38
rect -349 36 -347 38
rect -307 36 -305 38
rect -263 36 -261 38
rect -194 36 -192 38
rect -150 36 -148 38
rect -108 36 -106 38
rect -67 36 -65 38
rect -24 36 -22 38
rect 16 36 18 38
rect 59 36 61 38
rect -565 -27 -563 -25
rect -555 -27 -553 -25
rect -499 -20 -497 -18
rect -505 -30 -503 -28
rect -383 -27 -381 -25
rect -373 -27 -371 -25
rect -333 -27 -331 -25
rect -323 -27 -321 -25
rect -313 -27 -311 -25
rect -165 -27 -163 -25
rect -155 -27 -153 -25
rect -115 -27 -113 -25
rect -105 -27 -103 -25
rect -95 -27 -93 -25
rect -27 -27 -25 -25
rect -17 -27 -15 -25
rect 39 -20 41 -18
rect 33 -30 35 -28
rect -419 -107 -417 -105
rect -409 -107 -407 -105
rect -369 -107 -367 -105
rect -359 -107 -357 -105
rect -349 -107 -347 -105
rect -199 -107 -197 -105
rect -189 -107 -187 -105
rect -149 -107 -147 -105
rect -139 -107 -137 -105
rect -129 -107 -127 -105
rect -68 -107 -66 -105
rect -58 -107 -56 -105
rect -8 -104 -6 -102
rect -2 -114 0 -112
<< polyct1 >>
rect -516 44 -514 46
rect -526 36 -524 38
rect -476 44 -474 46
rect -486 36 -484 38
rect -433 44 -431 46
rect -443 36 -441 38
rect -329 44 -327 46
rect -339 36 -337 38
rect -287 44 -285 46
rect -297 36 -295 38
rect -243 44 -241 46
rect -253 36 -251 38
rect -174 44 -172 46
rect -184 36 -182 38
rect -130 44 -128 46
rect -140 36 -138 38
rect -88 44 -86 46
rect -98 36 -96 38
rect -47 44 -45 46
rect -57 36 -55 38
rect -4 44 -2 46
rect -14 36 -12 38
rect 36 44 38 46
rect 26 36 28 38
rect 79 44 81 46
rect 69 36 71 38
rect -545 -27 -543 -25
rect -538 -27 -536 -25
rect -519 -27 -517 -25
rect -472 -27 -470 -25
rect -448 -27 -446 -25
rect -422 -27 -420 -25
rect -408 -27 -406 -25
rect -343 -21 -341 -19
rect -295 -26 -293 -24
rect -347 -41 -345 -39
rect -254 -27 -252 -25
rect -230 -27 -228 -25
rect -204 -27 -202 -25
rect -190 -27 -188 -25
rect -125 -21 -123 -19
rect -77 -26 -75 -24
rect -272 -34 -270 -32
rect -129 -41 -127 -39
rect -7 -27 -5 -25
rect 0 -27 2 -25
rect 19 -27 21 -25
rect -54 -34 -52 -32
rect -383 -93 -381 -91
rect -508 -107 -506 -105
rect -484 -107 -482 -105
rect -458 -107 -456 -105
rect -444 -107 -442 -105
rect -331 -108 -329 -106
rect -379 -113 -377 -111
rect -308 -100 -306 -98
rect -163 -93 -161 -91
rect -288 -107 -286 -105
rect -264 -107 -262 -105
rect -238 -107 -236 -105
rect -224 -107 -222 -105
rect -111 -108 -109 -106
rect -159 -113 -157 -111
rect -88 -100 -86 -98
rect -48 -107 -46 -105
rect -41 -107 -39 -105
rect -22 -107 -20 -105
<< ndifct0 >>
rect -513 20 -511 22
rect -473 20 -471 22
rect -430 20 -428 22
rect -326 20 -324 22
rect -284 20 -282 22
rect -240 20 -238 22
rect -171 20 -169 22
rect -127 20 -125 22
rect -85 20 -83 22
rect -44 20 -42 22
rect -1 20 1 22
rect 39 20 41 22
rect 82 20 84 22
rect -559 -4 -557 -2
rect -542 -11 -540 -9
rect -532 -11 -530 -9
rect -532 -18 -530 -16
rect -522 -18 -520 -16
rect -512 -10 -510 -8
rect -502 -7 -500 -5
rect -455 -10 -453 -8
rect -465 -15 -463 -13
rect -416 -12 -414 -10
rect -406 -12 -404 -10
rect -351 -4 -349 -2
rect -362 -12 -360 -10
rect -340 -12 -338 -10
rect -310 -11 -308 -9
rect -300 -12 -298 -10
rect -290 -10 -288 -8
rect -237 -10 -235 -8
rect -279 -18 -277 -16
rect -247 -15 -245 -13
rect -198 -12 -196 -10
rect -188 -12 -186 -10
rect -133 -4 -131 -2
rect -144 -12 -142 -10
rect -122 -12 -120 -10
rect -92 -11 -90 -9
rect -82 -12 -80 -10
rect -72 -10 -70 -8
rect -21 -4 -19 -2
rect -61 -18 -59 -16
rect -4 -11 -2 -9
rect 6 -11 8 -9
rect 6 -18 8 -16
rect 16 -18 18 -16
rect 26 -10 28 -8
rect 36 -7 38 -5
rect -501 -119 -499 -117
rect -491 -124 -489 -122
rect -452 -122 -450 -120
rect -442 -122 -440 -120
rect -398 -122 -396 -120
rect -387 -130 -385 -128
rect -376 -122 -374 -120
rect -346 -123 -344 -121
rect -336 -122 -334 -120
rect -326 -124 -324 -122
rect -315 -116 -313 -114
rect -281 -119 -279 -117
rect -271 -124 -269 -122
rect -232 -122 -230 -120
rect -222 -122 -220 -120
rect -178 -122 -176 -120
rect -167 -130 -165 -128
rect -156 -122 -154 -120
rect -126 -123 -124 -121
rect -116 -122 -114 -120
rect -106 -124 -104 -122
rect -95 -116 -93 -114
rect -62 -130 -60 -128
rect -35 -116 -33 -114
rect -45 -123 -43 -121
rect -35 -123 -33 -121
rect -25 -116 -23 -114
rect -15 -124 -13 -122
rect -5 -127 -3 -125
<< ndifct1 >>
rect -543 22 -541 24
rect -503 22 -501 24
rect -460 22 -458 24
rect -532 10 -530 12
rect -356 22 -354 24
rect -492 10 -490 12
rect -314 22 -312 24
rect -449 10 -447 12
rect -270 22 -268 24
rect -345 10 -343 12
rect -201 22 -199 24
rect -303 10 -301 12
rect -157 22 -155 24
rect -259 10 -257 12
rect -115 22 -113 24
rect -190 10 -188 12
rect -74 22 -72 24
rect -146 10 -144 12
rect -31 22 -29 24
rect -104 10 -102 12
rect 9 22 11 24
rect -63 10 -61 12
rect 52 22 54 24
rect -20 10 -18 12
rect 20 10 22 12
rect 63 10 65 12
rect -570 -11 -568 -9
rect -444 -1 -442 1
rect -492 -11 -490 -9
rect -479 -18 -477 -16
rect -390 -1 -388 1
rect -426 -18 -424 -16
rect -372 -11 -370 -9
rect -328 -1 -326 1
rect -226 -1 -224 1
rect -261 -18 -259 -16
rect -172 -1 -170 1
rect -208 -18 -206 -16
rect -154 -11 -152 -9
rect -110 -1 -108 1
rect -32 -11 -30 -9
rect 46 -11 48 -9
rect -515 -116 -513 -114
rect -462 -116 -460 -114
rect -480 -133 -478 -131
rect -408 -123 -406 -121
rect -426 -133 -424 -131
rect -295 -116 -293 -114
rect -364 -133 -362 -131
rect -242 -116 -240 -114
rect -260 -133 -258 -131
rect -188 -123 -186 -121
rect -206 -133 -204 -131
rect -73 -123 -71 -121
rect -144 -133 -142 -131
rect 5 -123 7 -121
<< ntiect1 >>
rect -542 70 -540 72
rect -502 70 -500 72
rect -459 70 -457 72
rect -355 70 -353 72
rect -313 70 -311 72
rect -269 70 -267 72
rect -200 70 -198 72
rect -156 70 -154 72
rect -114 70 -112 72
rect -73 70 -71 72
rect -30 70 -28 72
rect 10 70 12 72
rect 53 70 55 72
rect -478 -61 -476 -59
rect -466 -61 -464 -59
rect -273 -61 -271 -59
rect -260 -61 -258 -59
rect -248 -61 -246 -59
rect -55 -61 -53 -59
rect -514 -73 -512 -71
rect -502 -73 -500 -71
rect -309 -73 -307 -71
rect -294 -73 -292 -71
rect -282 -73 -280 -71
rect -89 -73 -87 -71
<< ptiect1 >>
rect -542 10 -540 12
rect -502 10 -500 12
rect -459 10 -457 12
rect -355 10 -353 12
rect -313 10 -311 12
rect -269 10 -267 12
rect -200 10 -198 12
rect -156 10 -154 12
rect -114 10 -112 12
rect -73 10 -71 12
rect -30 10 -28 12
rect 10 10 12 12
rect 53 10 55 12
rect -478 -1 -476 1
rect -466 -1 -464 1
rect -273 -1 -271 1
rect -260 -1 -258 1
rect -248 -1 -246 1
rect -55 -1 -53 1
rect -514 -133 -512 -131
rect -502 -133 -500 -131
rect -309 -133 -307 -131
rect -294 -133 -292 -131
rect -282 -133 -280 -131
rect -89 -133 -87 -131
<< pdifct0 >>
rect -533 58 -531 60
rect -523 60 -521 62
rect -523 53 -521 55
rect -513 60 -511 62
rect -493 58 -491 60
rect -483 60 -481 62
rect -483 53 -481 55
rect -473 60 -471 62
rect -450 58 -448 60
rect -440 60 -438 62
rect -440 53 -438 55
rect -430 60 -428 62
rect -346 58 -344 60
rect -336 60 -334 62
rect -336 53 -334 55
rect -326 60 -324 62
rect -304 58 -302 60
rect -294 60 -292 62
rect -294 53 -292 55
rect -284 60 -282 62
rect -260 58 -258 60
rect -250 60 -248 62
rect -250 53 -248 55
rect -240 60 -238 62
rect -191 58 -189 60
rect -181 60 -179 62
rect -181 53 -179 55
rect -171 60 -169 62
rect -147 58 -145 60
rect -137 60 -135 62
rect -137 53 -135 55
rect -127 60 -125 62
rect -105 58 -103 60
rect -95 60 -93 62
rect -95 53 -93 55
rect -85 60 -83 62
rect -64 58 -62 60
rect -54 60 -52 62
rect -54 53 -52 55
rect -44 60 -42 62
rect -21 58 -19 60
rect -11 60 -9 62
rect -11 53 -9 55
rect -1 60 1 62
rect 19 58 21 60
rect 29 60 31 62
rect 29 53 31 55
rect 39 60 41 62
rect 62 58 64 60
rect 72 60 74 62
rect 72 53 74 55
rect 82 60 84 62
rect -560 -51 -558 -49
rect -560 -58 -558 -56
rect -550 -43 -548 -41
rect -550 -50 -548 -48
rect -538 -51 -536 -49
rect -538 -58 -536 -56
rect -515 -39 -513 -37
rect -503 -58 -501 -56
rect -468 -51 -466 -49
rect -452 -44 -450 -42
rect -452 -51 -450 -49
rect -442 -50 -440 -48
rect -442 -57 -440 -55
rect -415 -52 -413 -50
rect -405 -49 -403 -47
rect -390 -51 -388 -49
rect -405 -57 -403 -55
rect -370 -36 -368 -34
rect -370 -43 -368 -41
rect -360 -58 -358 -56
rect -350 -51 -348 -49
rect -340 -51 -338 -49
rect -330 -51 -328 -49
rect -340 -58 -338 -56
rect -320 -43 -318 -41
rect -310 -36 -308 -34
rect -310 -43 -308 -41
rect -289 -43 -287 -41
rect -279 -51 -277 -49
rect -300 -58 -298 -56
rect -250 -51 -248 -49
rect -234 -44 -232 -42
rect -234 -51 -232 -49
rect -224 -50 -222 -48
rect -224 -57 -222 -55
rect -197 -52 -195 -50
rect -187 -49 -185 -47
rect -172 -51 -170 -49
rect -187 -57 -185 -55
rect -152 -36 -150 -34
rect -152 -43 -150 -41
rect -142 -58 -140 -56
rect -132 -51 -130 -49
rect -122 -51 -120 -49
rect -112 -51 -110 -49
rect -122 -58 -120 -56
rect -102 -43 -100 -41
rect -92 -36 -90 -34
rect -92 -43 -90 -41
rect -71 -43 -69 -41
rect -61 -51 -59 -49
rect -82 -58 -80 -56
rect -22 -51 -20 -49
rect -22 -58 -20 -56
rect -12 -43 -10 -41
rect -12 -50 -10 -48
rect 0 -51 2 -49
rect 0 -58 2 -56
rect 23 -39 25 -37
rect 35 -58 37 -56
rect -504 -83 -502 -81
rect -488 -83 -486 -81
rect -488 -90 -486 -88
rect -478 -77 -476 -75
rect -478 -84 -476 -82
rect -451 -82 -449 -80
rect -441 -77 -439 -75
rect -441 -85 -439 -83
rect -426 -83 -424 -81
rect -406 -91 -404 -89
rect -406 -98 -404 -96
rect -396 -76 -394 -74
rect -386 -83 -384 -81
rect -376 -76 -374 -74
rect -376 -83 -374 -81
rect -366 -83 -364 -81
rect -356 -91 -354 -89
rect -346 -91 -344 -89
rect -346 -98 -344 -96
rect -336 -76 -334 -74
rect -325 -91 -323 -89
rect -315 -83 -313 -81
rect -284 -83 -282 -81
rect -268 -83 -266 -81
rect -268 -90 -266 -88
rect -258 -77 -256 -75
rect -258 -84 -256 -82
rect -231 -82 -229 -80
rect -221 -77 -219 -75
rect -221 -85 -219 -83
rect -206 -83 -204 -81
rect -186 -91 -184 -89
rect -186 -98 -184 -96
rect -176 -76 -174 -74
rect -166 -83 -164 -81
rect -156 -76 -154 -74
rect -156 -83 -154 -81
rect -146 -83 -144 -81
rect -136 -91 -134 -89
rect -126 -91 -124 -89
rect -126 -98 -124 -96
rect -116 -76 -114 -74
rect -105 -91 -103 -89
rect -95 -83 -93 -81
rect -63 -76 -61 -74
rect -63 -83 -61 -81
rect -53 -84 -51 -82
rect -53 -91 -51 -89
rect -41 -76 -39 -74
rect -41 -83 -39 -81
rect -6 -76 -4 -74
rect -18 -95 -16 -93
<< pdifct1 >>
rect -543 53 -541 55
rect -543 46 -541 48
rect -503 53 -501 55
rect -503 46 -501 48
rect -460 53 -458 55
rect -460 46 -458 48
rect -356 53 -354 55
rect -356 46 -354 48
rect -314 53 -312 55
rect -314 46 -312 48
rect -270 53 -268 55
rect -270 46 -268 48
rect -201 53 -199 55
rect -201 46 -199 48
rect -157 53 -155 55
rect -157 46 -155 48
rect -115 53 -113 55
rect -115 46 -113 48
rect -74 53 -72 55
rect -74 46 -72 48
rect -31 53 -29 55
rect -31 46 -29 48
rect 9 53 11 55
rect 9 46 11 48
rect 52 53 54 55
rect 52 46 54 48
rect -570 -36 -568 -34
rect -570 -43 -568 -41
rect -492 -39 -490 -37
rect -492 -46 -490 -44
rect -479 -36 -477 -34
rect -479 -43 -477 -41
rect -425 -36 -423 -34
rect -425 -43 -423 -41
rect -380 -43 -378 -41
rect -261 -36 -259 -34
rect -261 -43 -259 -41
rect -207 -36 -205 -34
rect -207 -43 -205 -41
rect -162 -43 -160 -41
rect -32 -36 -30 -34
rect -32 -43 -30 -41
rect 46 -39 48 -37
rect 46 -46 48 -44
rect -515 -91 -513 -89
rect -515 -98 -513 -96
rect -461 -91 -459 -89
rect -461 -98 -459 -96
rect -416 -91 -414 -89
rect -295 -91 -293 -89
rect -295 -98 -293 -96
rect -241 -91 -239 -89
rect -241 -98 -239 -96
rect -196 -91 -194 -89
rect -73 -91 -71 -89
rect -73 -98 -71 -96
rect 5 -88 7 -86
rect 5 -95 7 -93
<< alu0 >>
rect -535 60 -529 69
rect -535 58 -533 60
rect -531 58 -529 60
rect -535 57 -529 58
rect -524 62 -520 64
rect -524 60 -523 62
rect -521 60 -520 62
rect -524 55 -520 60
rect -515 62 -509 69
rect -515 60 -513 62
rect -511 60 -509 62
rect -515 59 -509 60
rect -495 60 -489 69
rect -495 58 -493 60
rect -491 58 -489 60
rect -495 57 -489 58
rect -484 62 -480 64
rect -484 60 -483 62
rect -481 60 -480 62
rect -524 54 -523 55
rect -537 53 -523 54
rect -521 53 -520 55
rect -537 50 -520 53
rect -537 38 -533 50
rect -484 55 -480 60
rect -475 62 -469 69
rect -475 60 -473 62
rect -471 60 -469 62
rect -475 59 -469 60
rect -452 60 -446 69
rect -452 58 -450 60
rect -448 58 -446 60
rect -452 57 -446 58
rect -441 62 -437 64
rect -441 60 -440 62
rect -438 60 -437 62
rect -484 54 -483 55
rect -497 53 -483 54
rect -481 53 -480 55
rect -497 50 -480 53
rect -537 36 -536 38
rect -534 36 -533 38
rect -537 31 -533 36
rect -537 27 -525 31
rect -541 24 -540 26
rect -529 23 -525 27
rect -497 38 -493 50
rect -441 55 -437 60
rect -432 62 -426 69
rect -432 60 -430 62
rect -428 60 -426 62
rect -432 59 -426 60
rect -348 60 -342 69
rect -348 58 -346 60
rect -344 58 -342 60
rect -348 57 -342 58
rect -337 62 -333 64
rect -337 60 -336 62
rect -334 60 -333 62
rect -441 54 -440 55
rect -454 53 -440 54
rect -438 53 -437 55
rect -454 50 -437 53
rect -497 36 -496 38
rect -494 36 -493 38
rect -497 31 -493 36
rect -497 27 -485 31
rect -501 24 -500 26
rect -529 22 -509 23
rect -529 20 -513 22
rect -511 20 -509 22
rect -529 19 -509 20
rect -489 23 -485 27
rect -454 38 -450 50
rect -337 55 -333 60
rect -328 62 -322 69
rect -328 60 -326 62
rect -324 60 -322 62
rect -328 59 -322 60
rect -306 60 -300 69
rect -306 58 -304 60
rect -302 58 -300 60
rect -306 57 -300 58
rect -295 62 -291 64
rect -295 60 -294 62
rect -292 60 -291 62
rect -337 54 -336 55
rect -350 53 -336 54
rect -334 53 -333 55
rect -350 50 -333 53
rect -454 36 -453 38
rect -451 36 -450 38
rect -454 31 -450 36
rect -454 27 -442 31
rect -458 24 -457 26
rect -489 22 -469 23
rect -489 20 -473 22
rect -471 20 -469 22
rect -489 19 -469 20
rect -446 23 -442 27
rect -350 38 -346 50
rect -295 55 -291 60
rect -286 62 -280 69
rect -286 60 -284 62
rect -282 60 -280 62
rect -286 59 -280 60
rect -262 60 -256 69
rect -262 58 -260 60
rect -258 58 -256 60
rect -262 57 -256 58
rect -251 62 -247 64
rect -251 60 -250 62
rect -248 60 -247 62
rect -295 54 -294 55
rect -308 53 -294 54
rect -292 53 -291 55
rect -308 50 -291 53
rect -350 36 -349 38
rect -347 36 -346 38
rect -350 31 -346 36
rect -350 27 -338 31
rect -354 24 -353 26
rect -446 22 -426 23
rect -446 20 -430 22
rect -428 20 -426 22
rect -446 19 -426 20
rect -342 23 -338 27
rect -308 38 -304 50
rect -251 55 -247 60
rect -242 62 -236 69
rect -242 60 -240 62
rect -238 60 -236 62
rect -242 59 -236 60
rect -193 60 -187 69
rect -193 58 -191 60
rect -189 58 -187 60
rect -193 57 -187 58
rect -182 62 -178 64
rect -182 60 -181 62
rect -179 60 -178 62
rect -251 54 -250 55
rect -264 53 -250 54
rect -248 53 -247 55
rect -264 50 -247 53
rect -308 36 -307 38
rect -305 36 -304 38
rect -308 31 -304 36
rect -308 27 -296 31
rect -312 24 -311 26
rect -342 22 -322 23
rect -342 20 -326 22
rect -324 20 -322 22
rect -342 19 -322 20
rect -300 23 -296 27
rect -264 38 -260 50
rect -182 55 -178 60
rect -173 62 -167 69
rect -173 60 -171 62
rect -169 60 -167 62
rect -173 59 -167 60
rect -149 60 -143 69
rect -149 58 -147 60
rect -145 58 -143 60
rect -149 57 -143 58
rect -138 62 -134 64
rect -138 60 -137 62
rect -135 60 -134 62
rect -182 54 -181 55
rect -195 53 -181 54
rect -179 53 -178 55
rect -195 50 -178 53
rect -264 36 -263 38
rect -261 36 -260 38
rect -264 31 -260 36
rect -264 27 -252 31
rect -268 24 -267 26
rect -300 22 -280 23
rect -300 20 -284 22
rect -282 20 -280 22
rect -300 19 -280 20
rect -256 23 -252 27
rect -195 38 -191 50
rect -138 55 -134 60
rect -129 62 -123 69
rect -129 60 -127 62
rect -125 60 -123 62
rect -129 59 -123 60
rect -107 60 -101 69
rect -107 58 -105 60
rect -103 58 -101 60
rect -107 57 -101 58
rect -96 62 -92 64
rect -96 60 -95 62
rect -93 60 -92 62
rect -138 54 -137 55
rect -151 53 -137 54
rect -135 53 -134 55
rect -151 50 -134 53
rect -195 36 -194 38
rect -192 36 -191 38
rect -195 31 -191 36
rect -195 27 -183 31
rect -199 24 -198 26
rect -256 22 -236 23
rect -256 20 -240 22
rect -238 20 -236 22
rect -256 19 -236 20
rect -187 23 -183 27
rect -151 38 -147 50
rect -96 55 -92 60
rect -87 62 -81 69
rect -87 60 -85 62
rect -83 60 -81 62
rect -87 59 -81 60
rect -66 60 -60 69
rect -66 58 -64 60
rect -62 58 -60 60
rect -66 57 -60 58
rect -55 62 -51 64
rect -55 60 -54 62
rect -52 60 -51 62
rect -96 54 -95 55
rect -109 53 -95 54
rect -93 53 -92 55
rect -109 50 -92 53
rect -151 36 -150 38
rect -148 36 -147 38
rect -151 31 -147 36
rect -151 27 -139 31
rect -155 24 -154 26
rect -187 22 -167 23
rect -187 20 -171 22
rect -169 20 -167 22
rect -187 19 -167 20
rect -143 23 -139 27
rect -109 38 -105 50
rect -55 55 -51 60
rect -46 62 -40 69
rect -46 60 -44 62
rect -42 60 -40 62
rect -46 59 -40 60
rect -23 60 -17 69
rect -23 58 -21 60
rect -19 58 -17 60
rect -23 57 -17 58
rect -12 62 -8 64
rect -12 60 -11 62
rect -9 60 -8 62
rect -55 54 -54 55
rect -68 53 -54 54
rect -52 53 -51 55
rect -68 50 -51 53
rect -109 36 -108 38
rect -106 36 -105 38
rect -109 31 -105 36
rect -109 27 -97 31
rect -113 24 -112 26
rect -143 22 -123 23
rect -143 20 -127 22
rect -125 20 -123 22
rect -143 19 -123 20
rect -101 23 -97 27
rect -68 38 -64 50
rect -12 55 -8 60
rect -3 62 3 69
rect -3 60 -1 62
rect 1 60 3 62
rect -3 59 3 60
rect 17 60 23 69
rect 17 58 19 60
rect 21 58 23 60
rect 17 57 23 58
rect 28 62 32 64
rect 28 60 29 62
rect 31 60 32 62
rect -12 54 -11 55
rect -25 53 -11 54
rect -9 53 -8 55
rect -25 50 -8 53
rect -68 36 -67 38
rect -65 36 -64 38
rect -68 31 -64 36
rect -68 27 -56 31
rect -72 24 -71 26
rect -101 22 -81 23
rect -101 20 -85 22
rect -83 20 -81 22
rect -101 19 -81 20
rect -60 23 -56 27
rect -25 38 -21 50
rect 28 55 32 60
rect 37 62 43 69
rect 37 60 39 62
rect 41 60 43 62
rect 37 59 43 60
rect 60 60 66 69
rect 60 58 62 60
rect 64 58 66 60
rect 60 57 66 58
rect 71 62 75 64
rect 71 60 72 62
rect 74 60 75 62
rect 28 54 29 55
rect 15 53 29 54
rect 31 53 32 55
rect 15 50 32 53
rect -25 36 -24 38
rect -22 36 -21 38
rect -25 31 -21 36
rect -25 27 -13 31
rect -29 24 -28 26
rect -60 22 -40 23
rect -60 20 -44 22
rect -42 20 -40 22
rect -60 19 -40 20
rect -17 23 -13 27
rect 15 38 19 50
rect 71 55 75 60
rect 80 62 86 69
rect 80 60 82 62
rect 84 60 86 62
rect 80 59 86 60
rect 71 54 72 55
rect 58 53 72 54
rect 74 53 75 55
rect 58 50 75 53
rect 15 36 16 38
rect 18 36 19 38
rect 15 31 19 36
rect 15 27 27 31
rect 11 24 12 26
rect -17 22 3 23
rect -17 20 -1 22
rect 1 20 3 22
rect -17 19 3 20
rect 23 23 27 27
rect 58 38 62 50
rect 58 36 59 38
rect 61 36 62 38
rect 58 31 62 36
rect 58 27 70 31
rect 54 24 55 26
rect 23 22 43 23
rect 23 20 39 22
rect 41 20 43 22
rect 23 19 43 20
rect 66 23 70 27
rect 66 22 86 23
rect 66 20 82 22
rect 84 20 86 22
rect 66 19 86 20
rect -561 -4 -559 -2
rect -557 -4 -555 -2
rect -561 -5 -555 -4
rect -503 -5 -499 -2
rect -503 -7 -502 -5
rect -500 -7 -499 -5
rect -533 -8 -508 -7
rect -548 -9 -538 -8
rect -548 -11 -542 -9
rect -540 -11 -538 -9
rect -548 -12 -538 -11
rect -533 -9 -512 -8
rect -533 -11 -532 -9
rect -530 -10 -512 -9
rect -510 -10 -508 -8
rect -503 -9 -499 -7
rect -530 -11 -508 -10
rect -548 -16 -544 -12
rect -564 -20 -544 -16
rect -564 -23 -560 -20
rect -566 -25 -560 -23
rect -566 -27 -565 -25
rect -563 -27 -560 -25
rect -566 -29 -560 -27
rect -564 -40 -560 -29
rect -556 -25 -552 -23
rect -533 -16 -529 -11
rect -533 -18 -532 -16
rect -530 -18 -529 -16
rect -533 -20 -529 -18
rect -524 -16 -509 -15
rect -524 -18 -522 -16
rect -520 -17 -509 -16
rect -520 -18 -495 -17
rect -524 -19 -499 -18
rect -513 -20 -499 -19
rect -497 -20 -495 -18
rect -513 -21 -495 -20
rect -556 -27 -555 -25
rect -553 -27 -552 -25
rect -556 -32 -552 -27
rect -513 -32 -509 -21
rect -516 -36 -509 -32
rect -506 -28 -502 -26
rect -506 -30 -505 -28
rect -503 -30 -502 -28
rect -516 -37 -512 -36
rect -516 -39 -515 -37
rect -513 -39 -512 -37
rect -564 -41 -524 -40
rect -516 -41 -512 -39
rect -506 -40 -502 -30
rect -564 -43 -550 -41
rect -548 -43 -524 -41
rect -564 -44 -524 -43
rect -508 -44 -502 -40
rect -551 -48 -547 -44
rect -528 -48 -504 -44
rect -466 -13 -462 -2
rect -457 -8 -412 -7
rect -457 -10 -455 -8
rect -453 -10 -412 -8
rect -457 -11 -416 -10
rect -418 -12 -416 -11
rect -414 -12 -412 -10
rect -418 -13 -412 -12
rect -408 -10 -402 -2
rect -353 -4 -351 -2
rect -349 -4 -347 -2
rect -353 -5 -347 -4
rect -291 -8 -287 -2
rect -408 -12 -406 -10
rect -404 -12 -402 -10
rect -408 -13 -402 -12
rect -363 -10 -359 -8
rect -332 -9 -306 -8
rect -363 -12 -362 -10
rect -360 -12 -359 -10
rect -477 -20 -476 -14
rect -466 -15 -465 -13
rect -463 -15 -462 -13
rect -466 -17 -462 -15
rect -477 -39 -476 -32
rect -453 -42 -431 -40
rect -453 -44 -452 -42
rect -450 -44 -431 -42
rect -562 -49 -556 -48
rect -562 -51 -560 -49
rect -558 -51 -556 -49
rect -562 -56 -556 -51
rect -551 -50 -550 -48
rect -548 -50 -547 -48
rect -551 -52 -547 -50
rect -540 -49 -534 -48
rect -540 -51 -538 -49
rect -536 -51 -534 -49
rect -562 -58 -560 -56
rect -558 -58 -556 -56
rect -540 -56 -534 -51
rect -470 -49 -464 -48
rect -470 -51 -468 -49
rect -466 -51 -464 -49
rect -540 -58 -538 -56
rect -536 -58 -534 -56
rect -505 -56 -499 -55
rect -505 -58 -503 -56
rect -501 -58 -499 -56
rect -470 -58 -464 -51
rect -453 -49 -449 -44
rect -453 -51 -452 -49
rect -450 -51 -449 -49
rect -453 -53 -449 -51
rect -444 -48 -438 -47
rect -444 -50 -442 -48
rect -440 -50 -438 -48
rect -444 -55 -438 -50
rect -435 -49 -431 -44
rect -363 -16 -359 -12
rect -384 -20 -359 -16
rect -353 -10 -336 -9
rect -353 -12 -340 -10
rect -338 -12 -336 -10
rect -353 -13 -336 -12
rect -332 -11 -310 -9
rect -308 -11 -306 -9
rect -332 -12 -306 -11
rect -301 -10 -297 -8
rect -301 -12 -300 -10
rect -298 -12 -297 -10
rect -291 -10 -290 -8
rect -288 -10 -287 -8
rect -291 -12 -287 -10
rect -384 -25 -380 -20
rect -353 -24 -349 -13
rect -384 -27 -383 -25
rect -381 -27 -380 -25
rect -384 -33 -380 -27
rect -375 -25 -349 -24
rect -375 -27 -373 -25
rect -371 -27 -349 -25
rect -375 -28 -349 -27
rect -332 -24 -328 -12
rect -301 -16 -297 -12
rect -280 -16 -276 -14
rect -384 -34 -366 -33
rect -384 -36 -370 -34
rect -368 -36 -366 -34
rect -384 -37 -366 -36
rect -372 -41 -366 -37
rect -372 -43 -370 -41
rect -368 -43 -366 -41
rect -372 -44 -366 -43
rect -406 -47 -402 -45
rect -406 -49 -405 -47
rect -403 -49 -402 -47
rect -362 -48 -358 -28
rect -335 -25 -328 -24
rect -335 -27 -333 -25
rect -331 -27 -328 -25
rect -335 -28 -328 -27
rect -332 -40 -328 -28
rect -324 -20 -297 -16
rect -324 -25 -320 -20
rect -324 -27 -323 -25
rect -321 -27 -320 -25
rect -324 -32 -320 -27
rect -315 -25 -300 -24
rect -315 -27 -313 -25
rect -311 -27 -300 -25
rect -315 -28 -300 -27
rect -324 -34 -307 -32
rect -324 -36 -310 -34
rect -308 -36 -307 -34
rect -332 -41 -316 -40
rect -332 -43 -320 -41
rect -318 -43 -316 -41
rect -332 -44 -316 -43
rect -311 -41 -307 -36
rect -311 -43 -310 -41
rect -308 -43 -307 -41
rect -311 -45 -307 -43
rect -304 -41 -300 -28
rect -280 -18 -279 -16
rect -277 -18 -276 -16
rect -280 -32 -276 -18
rect -248 -13 -244 -2
rect -239 -8 -194 -7
rect -239 -10 -237 -8
rect -235 -10 -194 -8
rect -239 -11 -198 -10
rect -200 -12 -198 -11
rect -196 -12 -194 -10
rect -200 -13 -194 -12
rect -190 -10 -184 -2
rect -135 -4 -133 -2
rect -131 -4 -129 -2
rect -135 -5 -129 -4
rect -73 -8 -69 -2
rect -23 -4 -21 -2
rect -19 -4 -17 -2
rect -23 -5 -17 -4
rect 35 -5 39 -2
rect 35 -7 36 -5
rect 38 -7 39 -5
rect 5 -8 30 -7
rect -190 -12 -188 -10
rect -186 -12 -184 -10
rect -190 -13 -184 -12
rect -145 -10 -141 -8
rect -114 -9 -88 -8
rect -145 -12 -144 -10
rect -142 -12 -141 -10
rect -290 -36 -276 -32
rect -290 -41 -286 -36
rect -304 -43 -289 -41
rect -287 -43 -286 -41
rect -304 -45 -286 -43
rect -259 -20 -258 -14
rect -248 -15 -247 -13
rect -245 -15 -244 -13
rect -248 -17 -244 -15
rect -259 -39 -258 -32
rect -235 -42 -213 -40
rect -235 -44 -234 -42
rect -232 -44 -213 -42
rect -304 -48 -300 -45
rect -435 -50 -411 -49
rect -435 -52 -415 -50
rect -413 -52 -411 -50
rect -435 -53 -411 -52
rect -444 -57 -442 -55
rect -440 -57 -438 -55
rect -444 -58 -438 -57
rect -406 -55 -402 -49
rect -392 -49 -346 -48
rect -392 -51 -390 -49
rect -388 -51 -350 -49
rect -348 -51 -346 -49
rect -392 -52 -346 -51
rect -342 -49 -336 -48
rect -342 -51 -340 -49
rect -338 -51 -336 -49
rect -406 -57 -405 -55
rect -403 -57 -402 -55
rect -406 -58 -402 -57
rect -362 -56 -356 -55
rect -362 -58 -360 -56
rect -358 -58 -356 -56
rect -342 -56 -336 -51
rect -332 -49 -300 -48
rect -332 -51 -330 -49
rect -328 -51 -300 -49
rect -332 -52 -300 -51
rect -281 -49 -275 -48
rect -281 -51 -279 -49
rect -277 -51 -275 -49
rect -342 -58 -340 -56
rect -338 -58 -336 -56
rect -302 -56 -296 -55
rect -302 -58 -300 -56
rect -298 -58 -296 -56
rect -281 -58 -275 -51
rect -252 -49 -246 -48
rect -252 -51 -250 -49
rect -248 -51 -246 -49
rect -252 -58 -246 -51
rect -235 -49 -231 -44
rect -235 -51 -234 -49
rect -232 -51 -231 -49
rect -235 -53 -231 -51
rect -226 -48 -220 -47
rect -226 -50 -224 -48
rect -222 -50 -220 -48
rect -226 -55 -220 -50
rect -217 -49 -213 -44
rect -145 -16 -141 -12
rect -166 -20 -141 -16
rect -135 -10 -118 -9
rect -135 -12 -122 -10
rect -120 -12 -118 -10
rect -135 -13 -118 -12
rect -114 -11 -92 -9
rect -90 -11 -88 -9
rect -114 -12 -88 -11
rect -83 -10 -79 -8
rect -83 -12 -82 -10
rect -80 -12 -79 -10
rect -73 -10 -72 -8
rect -70 -10 -69 -8
rect -73 -12 -69 -10
rect -10 -9 0 -8
rect -10 -11 -4 -9
rect -2 -11 0 -9
rect -10 -12 0 -11
rect 5 -9 26 -8
rect 5 -11 6 -9
rect 8 -10 26 -9
rect 28 -10 30 -8
rect 35 -9 39 -7
rect 8 -11 30 -10
rect -166 -25 -162 -20
rect -135 -24 -131 -13
rect -166 -27 -165 -25
rect -163 -27 -162 -25
rect -166 -33 -162 -27
rect -157 -25 -131 -24
rect -157 -27 -155 -25
rect -153 -27 -131 -25
rect -157 -28 -131 -27
rect -114 -24 -110 -12
rect -83 -16 -79 -12
rect -62 -16 -58 -14
rect -166 -34 -148 -33
rect -166 -36 -152 -34
rect -150 -36 -148 -34
rect -166 -37 -148 -36
rect -154 -41 -148 -37
rect -154 -43 -152 -41
rect -150 -43 -148 -41
rect -154 -44 -148 -43
rect -188 -47 -184 -45
rect -188 -49 -187 -47
rect -185 -49 -184 -47
rect -144 -48 -140 -28
rect -117 -25 -110 -24
rect -117 -27 -115 -25
rect -113 -27 -110 -25
rect -117 -28 -110 -27
rect -114 -40 -110 -28
rect -106 -20 -79 -16
rect -106 -25 -102 -20
rect -106 -27 -105 -25
rect -103 -27 -102 -25
rect -106 -32 -102 -27
rect -97 -25 -82 -24
rect -97 -27 -95 -25
rect -93 -27 -82 -25
rect -97 -28 -82 -27
rect -106 -34 -89 -32
rect -106 -36 -92 -34
rect -90 -36 -89 -34
rect -114 -41 -98 -40
rect -114 -43 -102 -41
rect -100 -43 -98 -41
rect -114 -44 -98 -43
rect -93 -41 -89 -36
rect -93 -43 -92 -41
rect -90 -43 -89 -41
rect -93 -45 -89 -43
rect -86 -41 -82 -28
rect -62 -18 -61 -16
rect -59 -18 -58 -16
rect -62 -32 -58 -18
rect -72 -36 -58 -32
rect -72 -41 -68 -36
rect -86 -43 -71 -41
rect -69 -43 -68 -41
rect -86 -45 -68 -43
rect -10 -16 -6 -12
rect -26 -20 -6 -16
rect -26 -23 -22 -20
rect -28 -25 -22 -23
rect -28 -27 -27 -25
rect -25 -27 -22 -25
rect -28 -29 -22 -27
rect -26 -40 -22 -29
rect -18 -25 -14 -23
rect 5 -16 9 -11
rect 5 -18 6 -16
rect 8 -18 9 -16
rect 5 -20 9 -18
rect 14 -16 29 -15
rect 14 -18 16 -16
rect 18 -17 29 -16
rect 18 -18 43 -17
rect 14 -19 39 -18
rect 25 -20 39 -19
rect 41 -20 43 -18
rect 25 -21 43 -20
rect -18 -27 -17 -25
rect -15 -27 -14 -25
rect -18 -32 -14 -27
rect 25 -32 29 -21
rect 22 -36 29 -32
rect 32 -28 36 -26
rect 32 -30 33 -28
rect 35 -30 36 -28
rect 22 -37 26 -36
rect 22 -39 23 -37
rect 25 -39 26 -37
rect -26 -41 14 -40
rect 22 -41 26 -39
rect 32 -40 36 -30
rect -26 -43 -12 -41
rect -10 -43 14 -41
rect -26 -44 14 -43
rect 30 -44 36 -40
rect -86 -48 -82 -45
rect -13 -48 -9 -44
rect 10 -48 34 -44
rect -217 -50 -193 -49
rect -217 -52 -197 -50
rect -195 -52 -193 -50
rect -217 -53 -193 -52
rect -226 -57 -224 -55
rect -222 -57 -220 -55
rect -226 -58 -220 -57
rect -188 -55 -184 -49
rect -174 -49 -128 -48
rect -174 -51 -172 -49
rect -170 -51 -132 -49
rect -130 -51 -128 -49
rect -174 -52 -128 -51
rect -124 -49 -118 -48
rect -124 -51 -122 -49
rect -120 -51 -118 -49
rect -188 -57 -187 -55
rect -185 -57 -184 -55
rect -188 -58 -184 -57
rect -144 -56 -138 -55
rect -144 -58 -142 -56
rect -140 -58 -138 -56
rect -124 -56 -118 -51
rect -114 -49 -82 -48
rect -114 -51 -112 -49
rect -110 -51 -82 -49
rect -114 -52 -82 -51
rect -63 -49 -57 -48
rect -63 -51 -61 -49
rect -59 -51 -57 -49
rect -124 -58 -122 -56
rect -120 -58 -118 -56
rect -84 -56 -78 -55
rect -84 -58 -82 -56
rect -80 -58 -78 -56
rect -63 -58 -57 -51
rect -24 -49 -18 -48
rect -24 -51 -22 -49
rect -20 -51 -18 -49
rect -24 -56 -18 -51
rect -13 -50 -12 -48
rect -10 -50 -9 -48
rect -13 -52 -9 -50
rect -2 -49 4 -48
rect -2 -51 0 -49
rect 2 -51 4 -49
rect -24 -58 -22 -56
rect -20 -58 -18 -56
rect -2 -56 4 -51
rect -2 -58 0 -56
rect 2 -58 4 -56
rect 33 -56 39 -55
rect 33 -58 35 -56
rect 37 -58 39 -56
rect -506 -81 -500 -74
rect -480 -75 -474 -74
rect -480 -77 -478 -75
rect -476 -77 -474 -75
rect -506 -83 -504 -81
rect -502 -83 -500 -81
rect -506 -84 -500 -83
rect -489 -81 -485 -79
rect -489 -83 -488 -81
rect -486 -83 -485 -81
rect -489 -88 -485 -83
rect -480 -82 -474 -77
rect -442 -75 -438 -74
rect -442 -77 -441 -75
rect -439 -77 -438 -75
rect -398 -76 -396 -74
rect -394 -76 -392 -74
rect -398 -77 -392 -76
rect -378 -76 -376 -74
rect -374 -76 -372 -74
rect -480 -84 -478 -82
rect -476 -84 -474 -82
rect -480 -85 -474 -84
rect -471 -80 -447 -79
rect -471 -82 -451 -80
rect -449 -82 -447 -80
rect -471 -83 -447 -82
rect -442 -83 -438 -77
rect -471 -88 -467 -83
rect -442 -85 -441 -83
rect -439 -85 -438 -83
rect -428 -81 -382 -80
rect -428 -83 -426 -81
rect -424 -83 -386 -81
rect -384 -83 -382 -81
rect -428 -84 -382 -83
rect -378 -81 -372 -76
rect -338 -76 -336 -74
rect -334 -76 -332 -74
rect -338 -77 -332 -76
rect -378 -83 -376 -81
rect -374 -83 -372 -81
rect -378 -84 -372 -83
rect -368 -81 -336 -80
rect -368 -83 -366 -81
rect -364 -83 -336 -81
rect -368 -84 -336 -83
rect -317 -81 -311 -74
rect -317 -83 -315 -81
rect -313 -83 -311 -81
rect -317 -84 -311 -83
rect -286 -81 -280 -74
rect -260 -75 -254 -74
rect -260 -77 -258 -75
rect -256 -77 -254 -75
rect -286 -83 -284 -81
rect -282 -83 -280 -81
rect -286 -84 -280 -83
rect -269 -81 -265 -79
rect -269 -83 -268 -81
rect -266 -83 -265 -81
rect -442 -87 -438 -85
rect -489 -90 -488 -88
rect -486 -90 -467 -88
rect -489 -92 -467 -90
rect -513 -100 -512 -93
rect -408 -89 -402 -88
rect -408 -91 -406 -89
rect -404 -91 -402 -89
rect -513 -118 -512 -112
rect -502 -117 -498 -115
rect -502 -119 -501 -117
rect -499 -119 -498 -117
rect -502 -130 -498 -119
rect -454 -120 -448 -119
rect -454 -121 -452 -120
rect -493 -122 -452 -121
rect -450 -122 -448 -120
rect -493 -124 -491 -122
rect -489 -124 -448 -122
rect -493 -125 -448 -124
rect -444 -120 -438 -119
rect -444 -122 -442 -120
rect -440 -122 -438 -120
rect -444 -130 -438 -122
rect -408 -95 -402 -91
rect -420 -96 -402 -95
rect -420 -98 -406 -96
rect -404 -98 -402 -96
rect -420 -99 -402 -98
rect -420 -105 -416 -99
rect -398 -104 -394 -84
rect -340 -87 -336 -84
rect -420 -107 -419 -105
rect -417 -107 -416 -105
rect -420 -112 -416 -107
rect -411 -105 -385 -104
rect -411 -107 -409 -105
rect -407 -107 -385 -105
rect -411 -108 -385 -107
rect -420 -116 -395 -112
rect -399 -120 -395 -116
rect -399 -122 -398 -120
rect -396 -122 -395 -120
rect -399 -124 -395 -122
rect -389 -119 -385 -108
rect -368 -89 -352 -88
rect -368 -91 -356 -89
rect -354 -91 -352 -89
rect -368 -92 -352 -91
rect -347 -89 -343 -87
rect -347 -91 -346 -89
rect -344 -91 -343 -89
rect -368 -104 -364 -92
rect -347 -96 -343 -91
rect -371 -105 -364 -104
rect -371 -107 -369 -105
rect -367 -107 -364 -105
rect -371 -108 -364 -107
rect -389 -120 -372 -119
rect -389 -122 -376 -120
rect -374 -122 -372 -120
rect -389 -123 -372 -122
rect -368 -120 -364 -108
rect -360 -98 -346 -96
rect -344 -98 -343 -96
rect -360 -100 -343 -98
rect -340 -89 -322 -87
rect -340 -91 -325 -89
rect -323 -91 -322 -89
rect -360 -105 -356 -100
rect -340 -104 -336 -91
rect -326 -96 -322 -91
rect -326 -100 -312 -96
rect -360 -107 -359 -105
rect -357 -107 -356 -105
rect -360 -112 -356 -107
rect -351 -105 -336 -104
rect -351 -107 -349 -105
rect -347 -107 -336 -105
rect -351 -108 -336 -107
rect -360 -116 -333 -112
rect -316 -114 -312 -100
rect -269 -88 -265 -83
rect -260 -82 -254 -77
rect -222 -75 -218 -74
rect -222 -77 -221 -75
rect -219 -77 -218 -75
rect -178 -76 -176 -74
rect -174 -76 -172 -74
rect -178 -77 -172 -76
rect -158 -76 -156 -74
rect -154 -76 -152 -74
rect -260 -84 -258 -82
rect -256 -84 -254 -82
rect -260 -85 -254 -84
rect -251 -80 -227 -79
rect -251 -82 -231 -80
rect -229 -82 -227 -80
rect -251 -83 -227 -82
rect -222 -83 -218 -77
rect -251 -88 -247 -83
rect -222 -85 -221 -83
rect -219 -85 -218 -83
rect -208 -81 -162 -80
rect -208 -83 -206 -81
rect -204 -83 -166 -81
rect -164 -83 -162 -81
rect -208 -84 -162 -83
rect -158 -81 -152 -76
rect -118 -76 -116 -74
rect -114 -76 -112 -74
rect -118 -77 -112 -76
rect -158 -83 -156 -81
rect -154 -83 -152 -81
rect -158 -84 -152 -83
rect -148 -81 -116 -80
rect -148 -83 -146 -81
rect -144 -83 -116 -81
rect -148 -84 -116 -83
rect -97 -81 -91 -74
rect -97 -83 -95 -81
rect -93 -83 -91 -81
rect -97 -84 -91 -83
rect -65 -76 -63 -74
rect -61 -76 -59 -74
rect -65 -81 -59 -76
rect -43 -76 -41 -74
rect -39 -76 -37 -74
rect -65 -83 -63 -81
rect -61 -83 -59 -81
rect -65 -84 -59 -83
rect -54 -82 -50 -80
rect -54 -84 -53 -82
rect -51 -84 -50 -82
rect -43 -81 -37 -76
rect -8 -76 -6 -74
rect -4 -76 -2 -74
rect -8 -77 -2 -76
rect -43 -83 -41 -81
rect -39 -83 -37 -81
rect -43 -84 -37 -83
rect -222 -87 -218 -85
rect -269 -90 -268 -88
rect -266 -90 -247 -88
rect -269 -92 -247 -90
rect -316 -116 -315 -114
rect -313 -116 -312 -114
rect -337 -120 -333 -116
rect -316 -118 -312 -116
rect -293 -100 -292 -93
rect -188 -89 -182 -88
rect -188 -91 -186 -89
rect -184 -91 -182 -89
rect -368 -121 -342 -120
rect -368 -123 -346 -121
rect -344 -123 -342 -121
rect -368 -124 -342 -123
rect -337 -122 -336 -120
rect -334 -122 -333 -120
rect -337 -124 -333 -122
rect -327 -122 -323 -120
rect -327 -124 -326 -122
rect -324 -124 -323 -122
rect -389 -128 -383 -127
rect -389 -130 -387 -128
rect -385 -130 -383 -128
rect -327 -130 -323 -124
rect -293 -118 -292 -112
rect -282 -117 -278 -115
rect -282 -119 -281 -117
rect -279 -119 -278 -117
rect -282 -130 -278 -119
rect -234 -120 -228 -119
rect -234 -121 -232 -120
rect -273 -122 -232 -121
rect -230 -122 -228 -120
rect -273 -124 -271 -122
rect -269 -124 -228 -122
rect -273 -125 -228 -124
rect -224 -120 -218 -119
rect -224 -122 -222 -120
rect -220 -122 -218 -120
rect -224 -130 -218 -122
rect -188 -95 -182 -91
rect -200 -96 -182 -95
rect -200 -98 -186 -96
rect -184 -98 -182 -96
rect -200 -99 -182 -98
rect -200 -105 -196 -99
rect -178 -104 -174 -84
rect -120 -87 -116 -84
rect -200 -107 -199 -105
rect -197 -107 -196 -105
rect -200 -112 -196 -107
rect -191 -105 -165 -104
rect -191 -107 -189 -105
rect -187 -107 -165 -105
rect -191 -108 -165 -107
rect -200 -116 -175 -112
rect -179 -120 -175 -116
rect -179 -122 -178 -120
rect -176 -122 -175 -120
rect -179 -124 -175 -122
rect -169 -119 -165 -108
rect -148 -89 -132 -88
rect -148 -91 -136 -89
rect -134 -91 -132 -89
rect -148 -92 -132 -91
rect -127 -89 -123 -87
rect -127 -91 -126 -89
rect -124 -91 -123 -89
rect -148 -104 -144 -92
rect -127 -96 -123 -91
rect -151 -105 -144 -104
rect -151 -107 -149 -105
rect -147 -107 -144 -105
rect -151 -108 -144 -107
rect -169 -120 -152 -119
rect -169 -122 -156 -120
rect -154 -122 -152 -120
rect -169 -123 -152 -122
rect -148 -120 -144 -108
rect -140 -98 -126 -96
rect -124 -98 -123 -96
rect -140 -100 -123 -98
rect -120 -89 -102 -87
rect -120 -91 -105 -89
rect -103 -91 -102 -89
rect -140 -105 -136 -100
rect -120 -104 -116 -91
rect -106 -96 -102 -91
rect -106 -100 -92 -96
rect -140 -107 -139 -105
rect -137 -107 -136 -105
rect -140 -112 -136 -107
rect -131 -105 -116 -104
rect -131 -107 -129 -105
rect -127 -107 -116 -105
rect -131 -108 -116 -107
rect -140 -116 -113 -112
rect -96 -114 -92 -100
rect -54 -88 -50 -84
rect -31 -88 -7 -84
rect -67 -89 -27 -88
rect -67 -91 -53 -89
rect -51 -91 -27 -89
rect -67 -92 -27 -91
rect -96 -116 -95 -114
rect -93 -116 -92 -114
rect -117 -120 -113 -116
rect -96 -118 -92 -116
rect -67 -103 -63 -92
rect -19 -93 -15 -91
rect -11 -92 -5 -88
rect -19 -95 -18 -93
rect -16 -95 -15 -93
rect -19 -96 -15 -95
rect -19 -100 -12 -96
rect -69 -105 -63 -103
rect -69 -107 -68 -105
rect -66 -107 -63 -105
rect -69 -109 -63 -107
rect -59 -105 -55 -100
rect -59 -107 -58 -105
rect -56 -107 -55 -105
rect -59 -109 -55 -107
rect -67 -112 -63 -109
rect -67 -116 -47 -112
rect -51 -120 -47 -116
rect -16 -111 -12 -100
rect -9 -102 -5 -92
rect -9 -104 -8 -102
rect -6 -104 -5 -102
rect -9 -106 -5 -104
rect -16 -112 2 -111
rect -36 -114 -32 -112
rect -16 -113 -2 -112
rect -36 -116 -35 -114
rect -33 -116 -32 -114
rect -148 -121 -122 -120
rect -148 -123 -126 -121
rect -124 -123 -122 -121
rect -148 -124 -122 -123
rect -117 -122 -116 -120
rect -114 -122 -113 -120
rect -117 -124 -113 -122
rect -107 -122 -103 -120
rect -107 -124 -106 -122
rect -104 -124 -103 -122
rect -51 -121 -41 -120
rect -51 -123 -45 -121
rect -43 -123 -41 -121
rect -51 -124 -41 -123
rect -36 -121 -32 -116
rect -27 -114 -2 -113
rect 0 -114 2 -112
rect -27 -116 -25 -114
rect -23 -115 2 -114
rect -23 -116 -12 -115
rect -27 -117 -12 -116
rect -36 -123 -35 -121
rect -33 -122 -11 -121
rect -33 -123 -15 -122
rect -36 -124 -15 -123
rect -13 -124 -11 -122
rect -169 -128 -163 -127
rect -169 -130 -167 -128
rect -165 -130 -163 -128
rect -107 -130 -103 -124
rect -36 -125 -11 -124
rect -6 -125 -2 -123
rect -6 -127 -5 -125
rect -3 -127 -2 -125
rect -64 -128 -58 -127
rect -64 -130 -62 -128
rect -60 -130 -58 -128
rect -6 -130 -2 -127
<< via1 >>
rect -512 53 -510 55
rect -472 53 -470 55
rect -520 35 -518 37
rect -539 19 -537 21
rect -480 36 -478 38
rect -503 19 -501 21
rect -429 48 -427 50
rect -460 19 -458 21
rect -436 27 -434 29
rect -325 48 -323 50
rect -283 53 -281 55
rect -353 19 -351 21
rect -333 28 -331 30
rect -239 53 -237 55
rect -291 36 -289 38
rect -315 19 -313 21
rect -271 28 -269 30
rect -170 53 -168 55
rect -247 28 -245 30
rect -126 53 -124 55
rect -199 19 -197 21
rect -178 28 -176 30
rect -150 20 -148 22
rect -134 28 -132 30
rect -84 48 -82 50
rect -43 52 -41 54
rect -92 36 -90 38
rect -116 19 -114 21
rect 0 53 2 55
rect -68 19 -66 21
rect -51 28 -49 30
rect -8 36 -6 38
rect -25 19 -23 21
rect 40 48 42 50
rect 83 53 85 55
rect 15 19 17 21
rect 33 27 35 29
rect 76 27 78 29
rect -539 -19 -537 -17
rect -523 -26 -521 -24
rect -472 -18 -470 -16
rect -440 -19 -438 -17
rect -407 -19 -405 -17
rect -448 -27 -446 -25
rect -472 -43 -470 -41
rect -500 -51 -498 -49
rect -416 -44 -414 -42
rect -343 -24 -341 -22
rect -387 -43 -385 -41
rect -295 -26 -293 -24
rect -271 -26 -269 -24
rect -279 -43 -277 -41
rect -254 -18 -252 -16
rect -222 -19 -220 -17
rect -199 -19 -197 -17
rect -189 -19 -187 -17
rect -230 -27 -228 -25
rect -254 -43 -252 -41
rect -198 -44 -196 -42
rect -125 -24 -123 -22
rect -166 -43 -164 -41
rect -77 -26 -75 -24
rect -53 -26 -51 -24
rect -61 -43 -59 -41
rect -1 -19 1 -17
rect -33 -39 -31 -37
rect 15 -26 17 -24
rect -452 -90 -450 -88
rect -484 -107 -482 -105
rect -508 -116 -506 -114
rect -476 -115 -474 -113
rect -443 -115 -441 -113
rect -379 -110 -377 -108
rect -315 -91 -313 -89
rect -331 -108 -329 -106
rect -232 -90 -230 -88
rect -264 -107 -262 -105
rect -288 -116 -286 -114
rect -241 -107 -239 -105
rect -256 -115 -254 -113
rect -223 -115 -221 -113
rect -159 -110 -157 -108
rect -95 -91 -93 -89
rect -111 -108 -109 -106
rect -34 -99 -32 -97
rect -51 -107 -49 -105
<< via2 >>
rect -472 68 -470 70
rect -512 57 -510 59
rect -239 68 -237 70
rect -283 57 -281 59
rect -170 57 -168 59
rect -126 57 -124 59
rect -43 58 -41 60
rect 0 58 2 60
rect 83 58 85 60
rect -429 44 -427 46
rect -325 44 -323 46
rect -84 44 -82 46
rect 40 44 42 46
rect -479 32 -477 34
rect -290 32 -288 34
rect -520 16 -518 18
rect -522 -12 -520 -10
rect -503 -12 -501 -10
rect -472 -13 -470 -11
rect -92 32 -90 34
rect -8 32 -6 34
rect -437 5 -435 7
rect -440 -13 -438 -11
rect -407 -15 -405 -13
rect -332 16 -330 18
rect -353 -15 -351 -13
rect -343 -17 -341 -15
rect -448 -35 -446 -33
rect -315 -35 -313 -33
rect -247 24 -245 26
rect -178 24 -176 26
rect -254 -13 -252 -11
rect -222 -13 -220 -11
rect -189 -15 -187 -13
rect -294 -35 -292 -33
rect -230 -35 -228 -33
rect -416 -50 -414 -48
rect -460 -61 -458 -59
rect -443 -61 -441 -59
rect -472 -84 -470 -82
rect -452 -84 -450 -82
rect -500 -99 -498 -97
rect -484 -99 -482 -97
rect -508 -121 -506 -119
rect -476 -121 -474 -119
rect -279 -50 -277 -48
rect -387 -63 -385 -61
rect -264 -63 -262 -61
rect -315 -84 -313 -82
rect -330 -99 -328 -97
rect -443 -119 -441 -117
rect -198 -50 -196 -48
rect -166 -61 -164 -59
rect -254 -84 -252 -82
rect -241 -84 -239 -82
rect -264 -99 -262 -97
rect -232 -84 -230 -82
rect -134 6 -132 8
rect -125 -17 -123 -15
rect 33 24 35 26
rect -50 16 -48 18
rect 76 24 78 26
rect -68 -11 -66 -9
rect -53 -11 -51 -9
rect -116 -35 -114 -33
rect -25 -11 -23 -9
rect -1 -11 1 -9
rect -76 -35 -74 -33
rect -61 -50 -59 -48
rect -51 -61 -49 -59
rect -150 -84 -148 -82
rect -95 -84 -93 -82
rect -110 -99 -108 -97
rect -379 -117 -377 -115
rect -288 -121 -286 -119
rect -256 -121 -254 -119
rect -223 -119 -221 -117
rect -159 -117 -157 -115
<< labels >>
rlabel alu1 25 9 25 9 6 vss
rlabel alu1 25 73 25 73 6 vdd
rlabel alu1 25 37 25 37 1 a0
rlabel alu1 33 33 33 33 1 a0
rlabel alu1 33 45 33 45 1 b1
rlabel alu1 41 53 41 53 1 b1
rlabel alu1 9 37 9 37 1 a0b1
rlabel alu1 17 21 17 21 1 a0b1
rlabel alu1 -15 9 -15 9 6 vss
rlabel alu1 -15 73 -15 73 6 vdd
rlabel alu1 -15 37 -15 37 1 a1
rlabel alu1 -7 33 -7 33 1 a1
rlabel alu1 -7 45 -7 45 1 b0
rlabel alu1 -31 37 -31 37 1 a1b0
rlabel alu1 -23 21 -23 21 1 a1b0
rlabel alu1 4 -62 4 -62 2 vdd
rlabel alu1 4 2 4 2 2 vss
rlabel ndifct1 -32 -10 -32 -10 1 c01
rlabel alu1 -24 -10 -24 -10 1 c01
rlabel alu1 -16 -10 -16 -10 1 c01
rlabel via1 -32 -38 -32 -38 1 c01
rlabel alu0 -5 -10 -5 -10 1 c01_inv
rlabel alu0 -24 -30 -24 -30 1 c01_inv
rlabel alu0 -11 -46 -11 -46 1 c01_inv
rlabel alu0 -6 -42 -6 -42 1 c01_inv
rlabel alu1 48 -26 48 -26 1 res1
rlabel alu1 40 -50 40 -50 1 res1
rlabel alu0 34 -35 34 -35 1 c01_inv
rlabel alu0 34 -19 34 -19 1 res1_inv
rlabel alu0 24 -36 24 -36 1 res1_inv
rlabel alu0 22 -17 22 -17 1 res1_inv
rlabel alu1 0 -22 0 -22 1 a1b0
rlabel alu1 -8 -26 -8 -26 1 a1b0
rlabel alu1 -16 -34 -16 -34 1 a0b1
rlabel alu1 -8 -34 -8 -34 1 a0b1
rlabel alu1 0 -34 0 -34 1 a0b1
rlabel alu1 8 -34 8 -34 1 a0b1
rlabel alu1 16 -30 16 -30 1 a0b1
rlabel alu1 68 9 68 9 6 vss
rlabel alu1 68 73 68 73 6 vdd
rlabel alu1 68 37 68 37 1 a0
rlabel alu1 76 33 76 33 1 a0
rlabel alu1 76 45 76 45 1 b0
rlabel alu1 1 53 1 53 1 b0
rlabel alu1 84 53 84 53 1 b0
rlabel alu1 52 37 52 37 1 res0
rlabel alu1 60 21 60 21 1 res0
rlabel alu0 76 21 76 21 1 res0_inv
rlabel alu0 60 40 60 40 1 res0_inv
rlabel alu1 -112 -62 -112 -62 8 vdd
rlabel alu1 -112 2 -112 2 8 vss
rlabel alu1 -209 -62 -209 -62 8 vdd
rlabel alu1 -209 2 -209 2 8 vss
rlabel alu1 -253 -62 -253 -62 8 vdd
rlabel alu1 -253 2 -253 2 8 vss
rlabel alu1 -261 -26 -261 -26 1 c02
rlabel via1 -253 -42 -253 -42 1 c02
rlabel alu1 -253 -22 -253 -22 1 c02_inv
rlabel alu1 -213 -18 -213 -18 1 c02_inv
rlabel alu1 -245 -26 -245 -26 1 c02_inv
rlabel alu1 -164 -42 -164 -42 1 s02
rlabel alu1 -172 -26 -172 -26 1 s02
rlabel alu1 -164 -10 -164 -10 1 s02
rlabel alu1 -156 -10 -156 -10 1 s02
rlabel alu0 -217 -9 -217 -9 1 fa_11_n3
rlabel alu0 -197 -10 -197 -10 1 fa_11_n3
rlabel alu0 -233 -46 -233 -46 1 fa_11_n1
rlabel alu0 -205 -51 -205 -51 1 fa_11_n1
rlabel alu1 -58 9 -58 9 6 vss
rlabel alu1 -58 73 -58 73 6 vdd
rlabel alu1 -58 37 -58 37 1 a2
rlabel alu1 -50 33 -50 33 1 a2
rlabel alu1 -50 45 -50 45 1 b0
rlabel via1 -42 53 -42 53 1 b0
rlabel alu1 -74 37 -74 37 1 a2b0
rlabel alu1 -66 21 -66 21 1 a2b0
rlabel polyct1 -52 -34 -52 -34 1 a2b0
rlabel alu1 -189 -30 -189 -30 1 a2b0
rlabel alu1 -99 73 -99 73 6 vdd
rlabel alu1 -99 9 -99 9 6 vss
rlabel alu1 -99 37 -99 37 1 a1
rlabel alu1 -91 33 -91 33 1 a1
rlabel alu1 -91 45 -91 45 1 b1
rlabel alu1 -83 53 -83 53 1 b1
rlabel alu1 -115 37 -115 37 1 a1b1
rlabel alu1 -237 -30 -237 -30 1 a1b1
rlabel alu1 -68 -22 -68 -22 1 a1b1
rlabel alu1 -107 21 -107 21 1 a1b1
rlabel alu1 -141 9 -141 9 6 vss
rlabel alu1 -141 73 -141 73 6 vdd
rlabel alu1 -141 37 -141 37 1 a3
rlabel alu1 -133 33 -133 33 1 a3
rlabel alu1 -125 53 -125 53 1 b0
rlabel alu1 -157 37 -157 37 1 a3b0
rlabel via1 -149 21 -149 21 1 a3b0
rlabel alu0 -149 40 -149 40 1 a3b0_inv
rlabel alu0 -136 57 -136 57 1 a3b0_inv
rlabel alu1 -133 45 -133 45 1 b0
rlabel alu1 -185 73 -185 73 6 vdd
rlabel alu1 -185 9 -185 9 6 vss
rlabel alu1 -177 45 -177 45 1 b2
rlabel alu1 -185 37 -185 37 1 a0
rlabel alu1 -177 33 -177 33 1 a0
rlabel alu1 -201 37 -201 37 1 a0b2
rlabel alu1 -193 21 -193 21 1 a0b2
rlabel alu1 -197 -18 -197 -18 1 a0b2
rlabel alu1 -205 -26 -205 -26 1 a0b2
rlabel alu1 -124 -30 -124 -30 1 a0b2
rlabel alu1 -132 -42 -132 -42 1 a0b2
rlabel alu0 -180 57 -180 57 1 a0b2_inv_0
rlabel alu0 -177 21 -177 21 1 a0b2_inv_0
rlabel alu0 -91 21 -91 21 1 a1b1_inv_0
rlabel alu0 -66 40 -66 40 1 a2b0_inv_0
rlabel alu0 -50 21 -50 21 1 a2b0_inv_0
rlabel alu0 -23 40 -23 40 1 a1b0_inv_0
rlabel alu0 -7 21 -7 21 1 a1b0_inv_0
rlabel alu0 17 40 17 40 1 a0b1_inv_0
rlabel alu0 33 21 33 21 1 a0b1_inv_0
rlabel alu0 -91 -38 -91 -38 1 a1b1_inv_1
rlabel alu0 -60 -25 -60 -25 1 a2b0_inv_1
rlabel alu0 -70 -38 -70 -38 1 a2b0_inv_1
rlabel alu0 -90 -26 -90 -26 1 a2b0_inv_1
rlabel alu0 -142 -38 -142 -38 1 a0b2_inv_1
rlabel alu0 -107 40 -107 40 1 a1b1_inv_0
rlabel alu1 -471 2 -471 2 8 vss
rlabel alu1 -471 -62 -471 -62 8 vdd
rlabel alu1 -427 2 -427 2 8 vss
rlabel alu1 -427 -62 -427 -62 8 vdd
rlabel alu1 -330 2 -330 2 8 vss
rlabel alu1 -330 -62 -330 -62 8 vdd
rlabel alu1 -479 -26 -479 -26 1 c03
rlabel via1 -471 -42 -471 -42 1 c03
rlabel alu1 -471 -22 -471 -22 1 c03_inv
rlabel alu1 -463 -26 -463 -26 1 c03_inv
rlabel alu1 -431 -18 -431 -18 1 c03_inv
rlabel alu1 -374 -10 -374 -10 1 s03
rlabel alu1 -382 -10 -382 -10 1 s03
rlabel alu1 -390 -26 -390 -26 1 s03
rlabel alu1 -382 -42 -382 -42 1 s03
rlabel alu0 -435 -9 -435 -9 1 fa_12_n3
rlabel alu0 -415 -10 -415 -10 1 fa_12_n3
rlabel alu0 -423 -51 -423 -51 1 fa_12_n1
rlabel alu0 -451 -46 -451 -46 1 fa_12_n1
rlabel alu1 -254 73 -254 73 6 vdd
rlabel alu1 -254 9 -254 9 6 vss
rlabel alu1 -238 53 -238 53 1 b3
rlabel alu1 -246 45 -246 45 1 b3
rlabel alu1 -254 37 -254 37 1 a0
rlabel alu1 -246 33 -246 33 1 a0
rlabel alu1 -270 37 -270 37 1 a0b3
rlabel alu1 -262 21 -262 21 1 a0b3
rlabel alu0 -249 57 -249 57 1 a0b3_inv_0
rlabel alu0 -262 40 -262 40 1 a0b3_inv_0
rlabel alu0 -246 21 -246 21 1 a0b3_inv_0
rlabel polyct1 -270 -34 -270 -34 1 a0b3
rlabel alu1 -415 -39 -415 -39 1 a0b3
rlabel alu1 -407 -30 -407 -30 1 a0b3
rlabel alu0 -278 -25 -278 -25 1 a0b3_inv_1
rlabel alu0 -288 -38 -288 -38 1 a0b3_inv_1
rlabel alu0 -308 -26 -308 -26 1 a0b3_inv_1
rlabel alu1 -298 73 -298 73 6 vdd
rlabel alu1 -298 9 -298 9 6 vss
rlabel alu1 -282 53 -282 53 1 b2
rlabel alu1 -290 45 -290 45 1 b2
rlabel alu1 -298 37 -298 37 1 a1
rlabel alu1 -290 33 -290 33 1 a1
rlabel alu1 -169 53 -169 53 1 b2
rlabel alu1 -314 37 -314 37 1 a1b2
rlabel alu1 -306 21 -306 21 1 a1b2
rlabel alu0 -293 57 -293 57 1 a1b2_inv_0
rlabel alu0 -306 40 -306 40 1 a1b2_inv_0
rlabel alu0 -290 21 -290 21 1 a1b2_inv_0
rlabel alu1 -286 -22 -286 -22 1 a1b2
rlabel alu1 -455 -30 -455 -30 1 a1b2
rlabel alu0 -299 -14 -299 -14 1 a1b2_inv_1
rlabel polyct0 -322 -26 -322 -26 1 a1b2_inv_1
rlabel alu0 -309 -38 -309 -38 1 a1b2_inv_1
rlabel alu1 -340 9 -340 9 6 vss
rlabel alu1 -340 73 -340 73 6 vdd
rlabel alu1 -324 53 -324 53 1 b1
rlabel alu1 -332 45 -332 45 1 b1
rlabel alu1 -340 37 -340 37 1 a2
rlabel alu1 -332 33 -332 33 1 a2
rlabel alu1 -356 37 -356 37 1 a2b1
rlabel alu0 -335 57 -335 57 1 a2b1_inv_0
rlabel alu0 -348 40 -348 40 1 a2b1_inv_0
rlabel alu1 -423 -26 -423 -26 1 a2b1
rlabel alu1 -415 -18 -415 -18 1 a2b1
rlabel alu1 -342 -30 -342 -30 1 a2b1
rlabel alu1 -350 -42 -350 -42 1 a2b1
rlabel alu0 -360 -38 -360 -38 1 a2b1_inv_1
rlabel alu0 -345 -11 -345 -11 1 a2b1_inv_1
rlabel alu1 -534 2 -534 2 2 vss
rlabel alu1 -534 -62 -534 -62 2 vdd
rlabel alu1 -570 -38 -570 -38 1 c04
rlabel ndifct1 -570 -10 -570 -10 1 c04
rlabel alu1 -562 -10 -562 -10 1 c04
rlabel alu1 -554 -10 -554 -10 1 c04
rlabel alu0 -562 -30 -562 -30 1 c04_inv_1
rlabel alu0 -544 -42 -544 -42 1 c04_inv_1
rlabel alu0 -549 -46 -549 -46 1 c04_inv_1
rlabel alu0 7 -13 7 -13 1 ha11
rlabel alu0 -504 -35 -504 -35 1 c04_inv_1
rlabel alu0 -543 -10 -543 -10 1 c04_inv_1
rlabel alu0 -531 -13 -531 -13 1 ha12
rlabel alu0 -520 -9 -520 -9 1 ha12
rlabel alu1 -490 -26 -490 -26 1 s04
rlabel alu1 -498 -50 -498 -50 1 s04
rlabel alu0 -516 -17 -516 -17 1 s04_inv_1
rlabel alu0 -504 -19 -504 -19 1 s04_inv_1
rlabel alu0 -514 -36 -514 -36 1 s04_inv_1
rlabel alu1 -348 21 -348 21 1 a2b1
rlabel alu1 -487 9 -487 9 6 vss
rlabel alu1 -487 73 -487 73 6 vdd
rlabel alu1 -527 9 -527 9 6 vss
rlabel alu1 -527 73 -527 73 6 vdd
rlabel alu1 -471 53 -471 53 1 b3
rlabel alu1 -479 45 -479 45 1 b3
rlabel alu1 -487 37 -487 37 1 a1
rlabel alu1 -479 33 -479 33 1 a1
rlabel alu1 -503 37 -503 37 1 a1b3
rlabel alu1 -495 21 -495 21 1 a1b3
rlabel alu0 -482 57 -482 57 1 a1b3_inv_0
rlabel alu0 -495 40 -495 40 1 a1b3_inv_0
rlabel alu0 -479 21 -479 21 1 a1b3_inv_0
rlabel alu1 -522 -30 -522 -30 1 a1b3
rlabel alu1 -530 -34 -530 -34 1 a1b3
rlabel alu1 -538 -34 -538 -34 1 a1b3
rlabel alu1 -546 -34 -546 -34 1 a1b3
rlabel alu1 -554 -34 -554 -34 1 a1b3
rlabel alu1 -527 37 -527 37 1 a2
rlabel alu1 -519 33 -519 33 1 a2
rlabel alu1 -519 45 -519 45 1 b2
rlabel alu1 -511 53 -511 53 1 b2
rlabel alu1 -543 37 -543 37 1 a2b2
rlabel alu0 -522 57 -522 57 1 a2b2_inv_0
rlabel alu0 -535 40 -535 40 1 a2b2_inv_0
rlabel alu0 -519 21 -519 21 1 a2b2_inv_0
rlabel alu1 -535 21 -535 21 1 a2b2
rlabel alu1 -538 -22 -538 -22 1 a2b2
rlabel alu1 -546 -26 -546 -26 1 a2b2
rlabel alu1 -37 -134 -37 -134 4 vss
rlabel alu1 -37 -70 -37 -70 4 vdd
rlabel alu1 -73 -94 -73 -94 1 c11
rlabel ndifct1 -73 -122 -73 -122 1 c11
rlabel alu1 -65 -122 -65 -122 1 c11
rlabel alu1 -57 -122 -57 -122 1 c11
rlabel alu0 -52 -86 -52 -86 1 c11_inv_2
rlabel alu0 -47 -90 -47 -90 1 c11_inv_2
rlabel alu0 -65 -102 -65 -102 1 c11_inv_2
rlabel alu0 -7 -97 -7 -97 1 c11_inv_2
rlabel alu1 7 -106 7 -106 1 res2
rlabel alu0 -7 -113 -7 -113 1 res2_inv
rlabel alu0 -19 -115 -19 -115 1 res2_inv
rlabel alu0 -34 -119 -34 -119 1 ha21
rlabel alu0 -23 -123 -23 -123 1 ha21
rlabel alu1 -57 -98 -57 -98 1 c01
rlabel alu1 -49 -98 -49 -98 1 c01
rlabel alu1 -41 -98 -41 -98 1 c01
rlabel alu1 -25 -102 -25 -102 1 c01
rlabel alu1 -41 -110 -41 -110 1 s02
rlabel alu0 -46 -122 -46 -122 1 c11_inv_2
rlabel alu0 -17 -96 -17 -96 1 res2_inv
rlabel alu1 -1 -82 -1 -82 1 res2
rlabel alu1 -287 -134 -287 -134 6 vss
rlabel alu1 -287 -70 -287 -70 6 vdd
rlabel alu1 -243 -134 -243 -134 6 vss
rlabel alu1 -243 -70 -243 -70 6 vdd
rlabel alu1 -146 -134 -146 -134 6 vss
rlabel alu1 -146 -70 -146 -70 6 vdd
rlabel alu1 -295 -106 -295 -106 1 c12
rlabel alu1 -287 -90 -287 -90 1 c12
rlabel alu1 -279 -106 -279 -106 1 c12_inv_2
rlabel alu1 -287 -110 -287 -110 1 c12_inv_2
rlabel alu1 -247 -114 -247 -114 1 c12_inv_2
rlabel alu0 -267 -86 -267 -86 1 fa_21_n1
rlabel alu0 -239 -81 -239 -81 1 fa_21_n1
rlabel alu0 -251 -123 -251 -123 1 fa_21_n3
rlabel alu0 -231 -122 -231 -122 1 fa_21_n3
rlabel alu1 -198 -90 -198 -90 1 s12
rlabel alu1 -206 -106 -206 -106 1 s12
rlabel alu1 -198 -122 -198 -122 1 s12
rlabel alu1 -190 -122 -190 -122 1 s12
rlabel alu1 -271 -102 -271 -102 1 s03
rlabel alu1 -102 -110 -102 -110 1 s03
rlabel polyct0 -138 -106 -138 -106 1 s03_inv_2
rlabel alu0 -115 -118 -115 -118 1 s03_inv_2
rlabel alu1 -86 -93 -86 -93 1 a3b0
rlabel alu1 -223 -102 -223 -102 1 a3b0
rlabel alu0 -124 -106 -124 -106 1 a3b0_inv_2
rlabel alu0 -104 -94 -104 -94 1 a3b0_inv_2
rlabel alu1 -231 -114 -231 -114 1 c02
rlabel alu1 -158 -102 -158 -102 1 c02
rlabel alu1 -166 -90 -166 -90 1 c02
rlabel alu0 -176 -94 -176 -94 1 c02_inv_2
rlabel alu0 -161 -121 -161 -121 1 c02_inv_2
rlabel alu0 -125 -94 -125 -94 1 s03_inv_2
rlabel alu0 -94 -107 -94 -107 1 a3b0_inv_2
rlabel alu1 -444 73 -444 73 6 vdd
rlabel alu1 -444 9 -444 9 6 vss
rlabel alu1 -444 37 -444 37 1 a3
rlabel alu0 -133 21 -133 21 1 a3b0_inv_0
rlabel alu1 -436 45 -436 45 1 b1
rlabel alu1 -428 53 -428 53 1 b1
rlabel alu1 -460 37 -460 37 1 a3b1
rlabel alu1 -452 21 -452 21 1 a3b1
rlabel alu0 -452 40 -452 40 1 a3b1_inv_0
rlabel alu1 -507 -134 -507 -134 6 vss
rlabel alu1 -507 -70 -507 -70 6 vdd
rlabel alu1 -463 -134 -463 -134 6 vss
rlabel alu1 -463 -70 -463 -70 6 vdd
rlabel alu1 -366 -134 -366 -134 6 vss
rlabel alu1 -366 -70 -366 -70 6 vdd
rlabel alu1 -507 -90 -507 -90 1 c13
rlabel alu1 -515 -106 -515 -106 1 c13
rlabel alu1 -499 -106 -499 -106 1 c13_inv_2
rlabel alu1 -507 -110 -507 -110 1 c13_inv_2
rlabel alu1 -467 -114 -467 -114 1 c13_inv_2
rlabel alu1 -426 -106 -426 -106 1 s13
rlabel alu1 -418 -90 -418 -90 1 s13
rlabel alu1 -418 -122 -418 -122 1 s13
rlabel alu1 -410 -122 -410 -122 1 s13
rlabel alu0 -459 -81 -459 -81 1 fa_22_n1
rlabel alu0 -487 -86 -487 -86 1 fa_22_n1
rlabel alu0 -471 -123 -471 -123 1 fa_22_n3
rlabel alu0 -451 -122 -451 -122 1 fa_22_n3
rlabel alu1 -491 -102 -491 -102 1 s04
rlabel alu1 -322 -110 -322 -110 1 s04
rlabel alu0 -335 -118 -335 -118 1 s04_inv_2
rlabel polyct0 -358 -106 -358 -106 1 s04_inv_2
rlabel alu0 -345 -94 -345 -94 1 s04_inv_2
rlabel alu1 -443 -102 -443 -102 1 c03
rlabel polyct1 -306 -98 -306 -98 1 c03
rlabel alu0 -314 -107 -314 -107 1 c03_inv_2
rlabel alu0 -324 -94 -324 -94 1 c03_inv_2
rlabel alu0 -344 -106 -344 -106 1 c03_inv_2
rlabel alu1 -451 -114 -451 -114 1 a3b1
rlabel alu1 -459 -106 -459 -106 1 a3b1
rlabel alu1 -378 -102 -378 -102 1 a3b1
rlabel alu1 -386 -90 -386 -90 1 a3b1
rlabel alu0 -396 -94 -396 -94 1 a3b1_inv_2
rlabel alu0 -381 -121 -381 -121 1 a3b1_inv_2
<< end >>
