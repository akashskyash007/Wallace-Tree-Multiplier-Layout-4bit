magic
tech scmos
timestamp 1684219586
<< ab >>
rect 58 -15 146 57
rect 147 -15 275 57
<< nwell >>
rect 53 17 280 62
<< pwell >>
rect 53 -20 280 17
<< poly >>
rect 94 50 96 55
rect 104 50 106 55
rect 111 50 113 55
rect 121 50 123 55
rect 131 50 133 55
rect 156 51 158 55
rect 166 51 168 55
rect 176 51 178 55
rect 186 51 188 55
rect 196 51 198 55
rect 216 51 218 55
rect 226 51 228 55
rect 236 51 238 55
rect 67 41 69 46
rect 186 34 188 37
rect 196 34 198 37
rect 186 32 198 34
rect 192 30 194 32
rect 196 30 198 32
rect 192 28 198 30
rect 247 44 249 48
rect 257 44 259 48
rect 247 27 249 30
rect 257 27 259 30
rect 247 25 273 27
rect 67 20 69 23
rect 94 20 96 23
rect 104 20 106 23
rect 67 18 73 20
rect 67 16 69 18
rect 71 16 73 18
rect 67 14 73 16
rect 91 18 106 20
rect 91 16 93 18
rect 95 16 106 18
rect 111 17 113 23
rect 121 20 123 23
rect 131 20 133 23
rect 156 20 158 23
rect 166 20 168 23
rect 176 20 178 23
rect 216 20 218 23
rect 226 20 228 23
rect 91 14 106 16
rect 110 14 113 17
rect 117 18 123 20
rect 117 16 119 18
rect 121 16 123 18
rect 117 14 123 16
rect 130 18 137 20
rect 130 16 133 18
rect 135 16 137 18
rect 130 14 137 16
rect 156 18 162 20
rect 156 16 158 18
rect 160 16 162 18
rect 156 14 162 16
rect 166 18 172 20
rect 176 18 212 20
rect 166 16 168 18
rect 170 16 172 18
rect 166 14 172 16
rect 67 11 69 14
rect 91 9 93 14
rect 103 11 105 14
rect 110 11 112 14
rect 120 11 122 14
rect 130 11 132 14
rect 67 -3 69 2
rect 157 5 159 14
rect 166 10 168 14
rect 184 10 186 18
rect 206 16 208 18
rect 210 16 212 18
rect 206 14 212 16
rect 216 18 222 20
rect 216 16 218 18
rect 220 16 222 18
rect 216 14 222 16
rect 226 18 232 20
rect 226 16 228 18
rect 230 16 232 18
rect 236 19 238 23
rect 236 17 250 19
rect 226 14 232 16
rect 244 15 246 17
rect 248 15 250 17
rect 196 12 202 14
rect 196 10 198 12
rect 200 10 202 12
rect 164 8 168 10
rect 164 5 166 8
rect 174 5 176 10
rect 91 -8 93 -3
rect 103 -6 105 -1
rect 110 -10 112 -1
rect 120 -6 122 -1
rect 130 -10 132 -1
rect 110 -12 132 -10
rect 196 8 202 10
rect 196 5 198 8
rect 219 5 221 14
rect 226 5 228 14
rect 244 13 250 15
rect 246 10 248 13
rect 257 11 259 25
rect 267 23 269 25
rect 271 23 273 25
rect 267 21 273 23
rect 236 5 238 10
rect 184 -7 186 -3
rect 157 -13 159 -8
rect 164 -13 166 -8
rect 174 -11 176 -8
rect 196 -11 198 -6
rect 174 -13 198 -11
rect 246 -7 248 -3
rect 219 -13 221 -8
rect 226 -13 228 -8
rect 236 -11 238 -8
rect 257 -11 259 0
rect 236 -13 259 -11
<< ndif >>
rect 60 9 67 11
rect 60 7 62 9
rect 64 7 67 9
rect 60 5 67 7
rect 62 2 67 5
rect 69 6 80 11
rect 95 9 103 11
rect 69 4 76 6
rect 78 4 80 6
rect 69 2 80 4
rect 86 3 91 9
rect 84 1 91 3
rect 84 -1 86 1
rect 88 -1 91 1
rect 84 -3 91 -1
rect 93 -1 103 9
rect 105 -1 110 11
rect 112 9 120 11
rect 112 7 115 9
rect 117 7 120 9
rect 112 -1 120 7
rect 122 3 130 11
rect 122 1 125 3
rect 127 1 130 3
rect 122 -1 130 1
rect 132 3 140 11
rect 179 5 184 10
rect 132 1 135 3
rect 137 1 140 3
rect 132 -1 140 1
rect 93 -3 101 -1
rect 95 -8 101 -3
rect 95 -10 97 -8
rect 99 -10 101 -8
rect 95 -12 101 -10
rect 149 -8 157 5
rect 159 -8 164 5
rect 166 2 174 5
rect 166 0 169 2
rect 171 0 174 2
rect 166 -8 174 0
rect 176 3 184 5
rect 176 1 179 3
rect 181 1 184 3
rect 176 -3 184 1
rect 186 5 194 10
rect 252 10 257 11
rect 241 5 246 10
rect 186 -3 196 5
rect 176 -8 181 -3
rect 188 -5 196 -3
rect 188 -7 190 -5
rect 192 -6 196 -5
rect 198 3 205 5
rect 198 1 201 3
rect 203 1 205 3
rect 198 -1 205 1
rect 198 -6 203 -1
rect 192 -7 194 -6
rect 149 -10 151 -8
rect 153 -10 155 -8
rect 149 -12 155 -10
rect 188 -9 194 -7
rect 211 -8 219 5
rect 221 -8 226 5
rect 228 2 236 5
rect 228 0 231 2
rect 233 0 236 2
rect 228 -8 236 0
rect 238 3 246 5
rect 238 1 241 3
rect 243 1 246 3
rect 238 -3 246 1
rect 248 1 257 10
rect 248 -1 251 1
rect 253 0 257 1
rect 259 9 266 11
rect 259 7 262 9
rect 264 7 266 9
rect 259 5 266 7
rect 259 0 264 5
rect 253 -1 255 0
rect 248 -3 255 -1
rect 238 -8 243 -3
rect 211 -10 213 -8
rect 215 -10 217 -8
rect 211 -12 217 -10
<< pdif >>
rect 89 44 94 50
rect 71 42 78 44
rect 71 41 73 42
rect 62 36 67 41
rect 60 34 67 36
rect 60 32 62 34
rect 64 32 67 34
rect 60 27 67 32
rect 60 25 62 27
rect 64 25 67 27
rect 60 23 67 25
rect 69 40 73 41
rect 75 40 78 42
rect 69 23 78 40
rect 87 42 94 44
rect 87 40 89 42
rect 91 40 94 42
rect 87 35 94 40
rect 87 33 89 35
rect 91 33 94 35
rect 87 31 94 33
rect 89 23 94 31
rect 96 48 104 50
rect 96 46 99 48
rect 101 46 104 48
rect 96 41 104 46
rect 96 39 99 41
rect 101 39 104 41
rect 96 23 104 39
rect 106 23 111 50
rect 113 34 121 50
rect 113 32 116 34
rect 118 32 121 34
rect 113 27 121 32
rect 113 25 116 27
rect 118 25 121 27
rect 113 23 121 25
rect 123 43 131 50
rect 123 41 126 43
rect 128 41 131 43
rect 123 23 131 41
rect 133 48 140 50
rect 133 46 136 48
rect 138 46 140 48
rect 133 40 140 46
rect 151 44 156 51
rect 133 38 136 40
rect 138 38 140 40
rect 149 42 156 44
rect 149 40 151 42
rect 153 40 156 42
rect 149 38 156 40
rect 133 23 140 38
rect 151 23 156 38
rect 158 34 166 51
rect 158 32 161 34
rect 163 32 166 34
rect 158 23 166 32
rect 168 34 176 51
rect 168 32 171 34
rect 173 32 176 34
rect 168 27 176 32
rect 168 25 171 27
rect 173 25 176 27
rect 168 23 176 25
rect 178 49 186 51
rect 178 47 181 49
rect 183 47 186 49
rect 178 37 186 47
rect 188 42 196 51
rect 188 40 191 42
rect 193 40 196 42
rect 188 37 196 40
rect 198 49 205 51
rect 198 47 201 49
rect 203 47 205 49
rect 198 42 205 47
rect 211 44 216 51
rect 198 40 201 42
rect 203 40 205 42
rect 198 37 205 40
rect 209 42 216 44
rect 209 40 211 42
rect 213 40 216 42
rect 209 38 216 40
rect 178 23 184 37
rect 211 23 216 38
rect 218 34 226 51
rect 218 32 221 34
rect 223 32 226 34
rect 218 23 226 32
rect 228 34 236 51
rect 228 32 231 34
rect 233 32 236 34
rect 228 27 236 32
rect 228 25 231 27
rect 233 25 236 27
rect 228 23 236 25
rect 238 49 245 51
rect 238 47 241 49
rect 243 47 245 49
rect 238 44 245 47
rect 238 30 247 44
rect 249 34 257 44
rect 249 32 252 34
rect 254 32 257 34
rect 249 30 257 32
rect 259 42 267 44
rect 259 40 262 42
rect 264 40 267 42
rect 259 30 267 40
rect 238 23 245 30
<< alu1 >>
rect 56 52 277 57
rect 56 50 63 52
rect 65 50 75 52
rect 77 50 268 52
rect 270 50 277 52
rect 56 49 277 50
rect 60 34 72 36
rect 60 32 62 34
rect 64 32 72 34
rect 60 30 72 32
rect 115 34 120 36
rect 115 32 116 34
rect 118 32 120 34
rect 60 27 64 30
rect 60 25 62 27
rect 60 9 64 25
rect 84 20 88 28
rect 115 27 120 32
rect 100 25 116 27
rect 118 25 120 27
rect 100 23 120 25
rect 124 35 128 36
rect 124 33 125 35
rect 127 33 128 35
rect 124 28 128 33
rect 149 34 165 35
rect 149 32 161 34
rect 163 32 165 34
rect 149 31 165 32
rect 124 23 137 28
rect 68 18 80 20
rect 68 16 69 18
rect 71 16 80 18
rect 68 14 80 16
rect 84 18 96 20
rect 84 16 93 18
rect 95 16 96 18
rect 84 14 96 16
rect 60 7 62 9
rect 60 -2 64 7
rect 68 9 72 14
rect 68 7 69 9
rect 71 7 72 9
rect 100 11 104 23
rect 115 18 127 19
rect 115 16 119 18
rect 121 16 127 18
rect 115 15 127 16
rect 131 18 137 23
rect 131 16 133 18
rect 135 16 137 18
rect 131 15 137 16
rect 123 11 127 15
rect 100 10 119 11
rect 100 8 101 10
rect 103 9 119 10
rect 103 8 115 9
rect 68 6 72 7
rect 100 7 115 8
rect 117 7 119 9
rect 123 10 137 11
rect 123 8 134 10
rect 136 8 137 10
rect 123 7 137 8
rect 100 6 119 7
rect 149 3 153 31
rect 188 32 201 35
rect 188 30 194 32
rect 196 30 201 32
rect 188 29 201 30
rect 149 2 173 3
rect 149 0 169 2
rect 171 0 173 2
rect 149 -1 173 0
rect 197 15 201 29
rect 197 13 198 15
rect 200 13 201 15
rect 197 12 201 13
rect 197 10 198 12
rect 200 10 201 12
rect 197 8 201 10
rect 260 34 273 36
rect 260 32 262 34
rect 264 32 273 34
rect 260 31 273 32
rect 269 27 273 31
rect 245 17 258 20
rect 245 15 246 17
rect 248 15 258 17
rect 245 14 258 15
rect 252 7 258 14
rect 268 25 273 27
rect 268 23 269 25
rect 271 23 273 25
rect 268 21 273 23
rect 269 14 273 21
rect 56 -8 277 -7
rect 56 -10 63 -8
rect 65 -10 75 -8
rect 77 -10 97 -8
rect 99 -10 151 -8
rect 153 -10 213 -8
rect 215 -10 268 -8
rect 270 -10 277 -8
rect 56 -15 277 -10
<< alu2 >>
rect 124 41 128 42
rect 124 39 125 41
rect 127 39 128 41
rect 124 35 128 39
rect 124 33 125 35
rect 127 33 128 35
rect 124 32 128 33
rect 261 41 265 42
rect 261 39 262 41
rect 264 39 265 41
rect 261 34 265 39
rect 261 32 262 34
rect 264 32 265 34
rect 261 31 265 32
rect 91 26 96 27
rect 91 24 93 26
rect 95 24 96 26
rect 91 18 96 24
rect 91 16 93 18
rect 95 16 96 18
rect 245 26 251 27
rect 245 24 247 26
rect 249 24 251 26
rect 245 17 251 24
rect 91 14 96 16
rect 197 15 201 16
rect 197 13 198 15
rect 200 13 201 15
rect 245 15 246 17
rect 248 15 251 17
rect 245 14 251 15
rect 100 10 104 11
rect 68 9 72 10
rect 68 7 69 9
rect 71 7 72 9
rect 68 4 72 7
rect 68 2 69 4
rect 71 2 72 4
rect 68 1 72 2
rect 100 8 101 10
rect 103 8 104 10
rect 100 4 104 8
rect 100 2 101 4
rect 103 2 104 4
rect 133 10 137 11
rect 133 8 134 10
rect 136 8 137 10
rect 133 6 137 8
rect 133 4 134 6
rect 136 4 137 6
rect 197 8 201 13
rect 197 6 198 8
rect 200 6 201 8
rect 197 4 201 6
rect 133 3 137 4
rect 100 1 104 2
<< alu3 >>
rect 124 41 265 42
rect 124 39 125 41
rect 127 39 262 41
rect 264 39 265 41
rect 124 38 265 39
rect 91 26 251 27
rect 91 24 93 26
rect 95 24 247 26
rect 249 24 251 26
rect 91 23 251 24
rect 197 8 201 9
rect 197 7 198 8
rect 133 6 198 7
rect 200 6 201 8
rect 68 4 105 5
rect 68 2 69 4
rect 71 2 101 4
rect 103 2 105 4
rect 133 4 134 6
rect 136 4 201 6
rect 133 3 201 4
rect 68 1 105 2
<< ptie >>
rect 61 -8 79 -6
rect 61 -10 63 -8
rect 65 -10 75 -8
rect 77 -10 79 -8
rect 61 -12 79 -10
rect 266 -8 272 -6
rect 266 -10 268 -8
rect 270 -10 272 -8
rect 266 -12 272 -10
<< ntie >>
rect 61 52 79 54
rect 61 50 63 52
rect 65 50 75 52
rect 77 50 79 52
rect 266 52 272 54
rect 61 48 79 50
rect 266 50 268 52
rect 270 50 272 52
rect 266 48 272 50
<< nmos >>
rect 67 2 69 11
rect 91 -3 93 9
rect 103 -1 105 11
rect 110 -1 112 11
rect 120 -1 122 11
rect 130 -1 132 11
rect 157 -8 159 5
rect 164 -8 166 5
rect 174 -8 176 5
rect 184 -3 186 10
rect 196 -6 198 5
rect 219 -8 221 5
rect 226 -8 228 5
rect 236 -8 238 5
rect 246 -3 248 10
rect 257 0 259 11
<< pmos >>
rect 67 23 69 41
rect 94 23 96 50
rect 104 23 106 50
rect 111 23 113 50
rect 121 23 123 50
rect 131 23 133 50
rect 156 23 158 51
rect 166 23 168 51
rect 176 23 178 51
rect 186 37 188 51
rect 196 37 198 51
rect 216 23 218 51
rect 226 23 228 51
rect 236 23 238 51
rect 247 30 249 44
rect 257 30 259 44
<< polyct0 >>
rect 158 16 160 18
rect 168 16 170 18
rect 208 16 210 18
rect 218 16 220 18
rect 228 16 230 18
<< polyct1 >>
rect 194 30 196 32
rect 69 16 71 18
rect 93 16 95 18
rect 119 16 121 18
rect 133 16 135 18
rect 246 15 248 17
rect 198 10 200 12
rect 269 23 271 25
<< ndifct0 >>
rect 76 4 78 6
rect 86 -1 88 1
rect 125 1 127 3
rect 135 1 137 3
rect 179 1 181 3
rect 190 -7 192 -5
rect 201 1 203 3
rect 231 0 233 2
rect 241 1 243 3
rect 251 -1 253 1
rect 262 7 264 9
<< ndifct1 >>
rect 62 7 64 9
rect 115 7 117 9
rect 97 -10 99 -8
rect 169 0 171 2
rect 151 -10 153 -8
rect 213 -10 215 -8
<< ntiect1 >>
rect 63 50 65 52
rect 75 50 77 52
rect 268 50 270 52
<< ptiect1 >>
rect 63 -10 65 -8
rect 75 -10 77 -8
rect 268 -10 270 -8
<< pdifct0 >>
rect 73 40 75 42
rect 89 40 91 42
rect 89 33 91 35
rect 99 46 101 48
rect 99 39 101 41
rect 126 41 128 43
rect 136 46 138 48
rect 136 38 138 40
rect 151 40 153 42
rect 171 32 173 34
rect 171 25 173 27
rect 181 47 183 49
rect 191 40 193 42
rect 201 47 203 49
rect 201 40 203 42
rect 211 40 213 42
rect 221 32 223 34
rect 231 32 233 34
rect 231 25 233 27
rect 241 47 243 49
rect 252 32 254 34
rect 262 40 264 42
<< pdifct1 >>
rect 62 32 64 34
rect 62 25 64 27
rect 116 32 118 34
rect 116 25 118 27
rect 161 32 163 34
<< alu0 >>
rect 71 42 77 49
rect 97 48 103 49
rect 97 46 99 48
rect 101 46 103 48
rect 71 40 73 42
rect 75 40 77 42
rect 71 39 77 40
rect 88 42 92 44
rect 88 40 89 42
rect 91 40 92 42
rect 88 35 92 40
rect 97 41 103 46
rect 135 48 139 49
rect 135 46 136 48
rect 138 46 139 48
rect 179 47 181 49
rect 183 47 185 49
rect 179 46 185 47
rect 199 47 201 49
rect 203 47 205 49
rect 97 39 99 41
rect 101 39 103 41
rect 97 38 103 39
rect 106 43 130 44
rect 106 41 126 43
rect 128 41 130 43
rect 106 40 130 41
rect 135 40 139 46
rect 106 35 110 40
rect 135 38 136 40
rect 138 38 139 40
rect 149 42 195 43
rect 149 40 151 42
rect 153 40 191 42
rect 193 40 195 42
rect 149 39 195 40
rect 199 42 205 47
rect 239 47 241 49
rect 243 47 245 49
rect 239 46 245 47
rect 199 40 201 42
rect 203 40 205 42
rect 199 39 205 40
rect 209 42 241 43
rect 209 40 211 42
rect 213 40 241 42
rect 209 39 241 40
rect 260 42 266 49
rect 260 40 262 42
rect 264 40 266 42
rect 260 39 266 40
rect 135 36 139 38
rect 88 33 89 35
rect 91 33 110 35
rect 88 31 110 33
rect 64 23 65 30
rect 169 34 175 35
rect 169 32 171 34
rect 173 32 175 34
rect 64 5 65 11
rect 75 6 79 8
rect 75 4 76 6
rect 78 4 79 6
rect 75 -7 79 4
rect 123 3 129 4
rect 123 2 125 3
rect 84 1 125 2
rect 127 1 129 3
rect 84 -1 86 1
rect 88 -1 129 1
rect 84 -2 129 -1
rect 133 3 139 4
rect 133 1 135 3
rect 137 1 139 3
rect 133 -7 139 1
rect 169 28 175 32
rect 157 27 175 28
rect 157 25 171 27
rect 173 25 175 27
rect 157 24 175 25
rect 157 18 161 24
rect 179 19 183 39
rect 237 36 241 39
rect 157 16 158 18
rect 160 16 161 18
rect 157 11 161 16
rect 166 18 192 19
rect 166 16 168 18
rect 170 16 192 18
rect 166 15 192 16
rect 157 7 182 11
rect 178 3 182 7
rect 178 1 179 3
rect 181 1 182 3
rect 178 -1 182 1
rect 188 4 192 15
rect 209 34 225 35
rect 209 32 221 34
rect 223 32 225 34
rect 209 31 225 32
rect 230 34 234 36
rect 230 32 231 34
rect 233 32 234 34
rect 209 19 213 31
rect 230 27 234 32
rect 206 18 213 19
rect 206 16 208 18
rect 210 16 213 18
rect 206 15 213 16
rect 188 3 205 4
rect 188 1 201 3
rect 203 1 205 3
rect 188 0 205 1
rect 209 3 213 15
rect 217 25 231 27
rect 233 25 234 27
rect 217 23 234 25
rect 237 34 255 36
rect 237 32 252 34
rect 254 32 255 34
rect 217 18 221 23
rect 237 19 241 32
rect 251 27 255 32
rect 251 23 265 27
rect 217 16 218 18
rect 220 16 221 18
rect 217 11 221 16
rect 226 18 241 19
rect 226 16 228 18
rect 230 16 241 18
rect 226 15 241 16
rect 217 7 244 11
rect 261 9 265 23
rect 261 7 262 9
rect 264 7 265 9
rect 240 3 244 7
rect 261 5 265 7
rect 209 2 235 3
rect 209 0 231 2
rect 233 0 235 2
rect 209 -1 235 0
rect 240 1 241 3
rect 243 1 244 3
rect 240 -1 244 1
rect 250 1 254 3
rect 250 -1 251 1
rect 253 -1 254 1
rect 188 -5 194 -4
rect 188 -7 190 -5
rect 192 -7 194 -5
rect 250 -7 254 -1
<< via1 >>
rect 125 33 127 35
rect 93 16 95 18
rect 69 7 71 9
rect 101 8 103 10
rect 134 8 136 10
rect 198 13 200 15
rect 262 32 264 34
rect 246 15 248 17
<< via2 >>
rect 125 39 127 41
rect 262 39 264 41
rect 93 24 95 26
rect 247 24 249 26
rect 69 2 71 4
rect 101 2 103 4
rect 134 4 136 6
rect 198 6 200 8
<< labels >>
rlabel via1 263 33 263 33 6 b
rlabel alu1 271 25 271 25 6 b
rlabel alu1 255 13 255 13 6 a
rlabel alu1 247 17 247 17 6 a
rlabel alu1 211 53 211 53 6 vdd
rlabel alu1 211 -11 211 -11 6 vss
rlabel alu1 191 33 191 33 6 c
rlabel alu1 199 21 199 21 6 c
rlabel alu0 225 41 225 41 6 bn
rlabel alu0 263 16 263 16 6 bn
rlabel alu0 253 29 253 29 6 bn
rlabel alu0 233 17 233 17 6 bn
rlabel alu0 242 5 242 5 6 an
rlabel polyct0 219 17 219 17 6 an
rlabel alu0 232 29 232 29 6 an
rlabel alu0 181 29 181 29 6 cn
rlabel alu0 172 41 172 41 6 cn
rlabel alu0 196 2 196 2 6 cn
rlabel alu1 134 21 134 21 6 b
rlabel alu1 134 9 134 9 6 c
rlabel alu1 114 53 114 53 6 vdd
rlabel alu1 126 33 126 33 6 b
rlabel alu1 126 9 126 9 6 c
rlabel alu1 118 17 118 17 6 c
rlabel alu1 114 -11 114 -11 6 vss
rlabel alu1 86 21 86 21 6 a
rlabel polyct1 94 17 94 17 6 a
rlabel alu0 118 42 118 42 6 n1
rlabel alu0 126 1 126 1 6 n3
rlabel alu0 106 0 106 0 6 n3
rlabel alu0 90 37 90 37 6 n1
rlabel alu1 70 53 70 53 6 vdd
rlabel alu1 70 -11 70 -11 6 vss
rlabel alu1 78 17 78 17 1 cout_inv
rlabel alu1 70 13 70 13 1 cout_inv
rlabel alu1 62 17 62 17 1 cout
rlabel alu1 70 33 70 33 1 cout
rlabel alu1 110 9 110 9 1 cout_inv
rlabel alu1 159 33 159 33 1 sum
rlabel alu1 151 17 151 17 1 sum
rlabel alu1 159 1 159 1 1 sum
rlabel alu1 167 1 167 1 1 sum
<< end >>
