magic
tech scmos
timestamp 1684940948
<< ab >>
rect 40 149 120 220
rect 123 149 163 220
rect 227 149 267 220
rect 269 149 309 220
rect 313 149 353 220
rect 382 149 422 220
rect 426 149 466 220
rect 468 149 508 220
rect 509 149 549 220
rect 552 149 632 220
rect 635 149 675 220
rect -77 77 -37 149
rect -35 148 192 149
rect -35 77 101 148
rect 104 77 192 148
rect 193 148 675 149
rect 193 77 321 148
rect 322 77 410 148
rect 411 77 539 148
rect 543 77 639 148
rect -194 5 -154 77
rect -150 5 -62 77
rect -61 5 67 77
rect 68 5 156 77
rect 157 5 285 77
rect 288 5 376 77
rect 377 5 598 77
rect -212 -67 -124 5
rect -123 -67 5 5
rect 8 -67 96 5
rect 97 -67 313 5
rect 314 -67 442 5
rect 445 -67 541 5
<< nwell >>
rect 35 180 680 225
rect -82 82 644 117
rect -199 72 644 82
rect -199 37 603 72
rect -217 -72 546 -27
<< pwell >>
rect 35 154 680 180
rect -82 143 680 154
rect -82 117 644 143
rect -199 10 603 37
rect -217 0 603 10
rect -217 -27 546 0
<< poly >>
rect 49 205 51 209
rect 59 207 61 212
rect 69 207 71 212
rect 89 205 91 209
rect 99 207 101 212
rect 109 207 111 212
rect 49 183 51 187
rect 59 183 61 194
rect 69 191 71 194
rect 69 189 75 191
rect 69 187 71 189
rect 73 187 75 189
rect 132 205 134 209
rect 142 207 144 212
rect 152 207 154 212
rect 69 185 75 187
rect 49 181 55 183
rect 49 179 51 181
rect 53 179 55 181
rect 49 177 55 179
rect 59 181 65 183
rect 59 179 61 181
rect 63 179 65 181
rect 59 177 65 179
rect 49 172 51 177
rect 62 172 64 177
rect 69 172 71 185
rect 89 183 91 187
rect 99 183 101 194
rect 109 191 111 194
rect 109 189 115 191
rect 109 187 111 189
rect 113 187 115 189
rect 236 205 238 209
rect 246 207 248 212
rect 256 207 258 212
rect 109 185 115 187
rect 89 181 95 183
rect 89 179 91 181
rect 93 179 95 181
rect 89 177 95 179
rect 99 181 105 183
rect 99 179 101 181
rect 103 179 105 181
rect 99 177 105 179
rect 89 172 91 177
rect 102 172 104 177
rect 109 172 111 185
rect 132 183 134 187
rect 142 183 144 194
rect 152 191 154 194
rect 152 189 158 191
rect 152 187 154 189
rect 156 187 158 189
rect 278 205 280 209
rect 288 207 290 212
rect 298 207 300 212
rect 152 185 158 187
rect 132 181 138 183
rect 132 179 134 181
rect 136 179 138 181
rect 132 177 138 179
rect 142 181 148 183
rect 142 179 144 181
rect 146 179 148 181
rect 142 177 148 179
rect 132 172 134 177
rect 145 172 147 177
rect 152 172 154 185
rect 236 183 238 187
rect 246 183 248 194
rect 256 191 258 194
rect 256 189 262 191
rect 256 187 258 189
rect 260 187 262 189
rect 322 205 324 209
rect 332 207 334 212
rect 342 207 344 212
rect 256 185 262 187
rect 236 181 242 183
rect 236 179 238 181
rect 240 179 242 181
rect 236 177 242 179
rect 246 181 252 183
rect 246 179 248 181
rect 250 179 252 181
rect 246 177 252 179
rect 236 172 238 177
rect 249 172 251 177
rect 256 172 258 185
rect 278 183 280 187
rect 288 183 290 194
rect 298 191 300 194
rect 298 189 304 191
rect 298 187 300 189
rect 302 187 304 189
rect 391 205 393 209
rect 401 207 403 212
rect 411 207 413 212
rect 298 185 304 187
rect 278 181 284 183
rect 278 179 280 181
rect 282 179 284 181
rect 278 177 284 179
rect 288 181 294 183
rect 288 179 290 181
rect 292 179 294 181
rect 288 177 294 179
rect 278 172 280 177
rect 291 172 293 177
rect 298 172 300 185
rect 322 183 324 187
rect 332 183 334 194
rect 342 191 344 194
rect 342 189 348 191
rect 342 187 344 189
rect 346 187 348 189
rect 435 205 437 209
rect 445 207 447 212
rect 455 207 457 212
rect 342 185 348 187
rect 322 181 328 183
rect 322 179 324 181
rect 326 179 328 181
rect 322 177 328 179
rect 332 181 338 183
rect 332 179 334 181
rect 336 179 338 181
rect 332 177 338 179
rect 322 172 324 177
rect 335 172 337 177
rect 342 172 344 185
rect 391 183 393 187
rect 401 183 403 194
rect 411 191 413 194
rect 411 189 417 191
rect 411 187 413 189
rect 415 187 417 189
rect 477 205 479 209
rect 487 207 489 212
rect 497 207 499 212
rect 411 185 417 187
rect 391 181 397 183
rect 391 179 393 181
rect 395 179 397 181
rect 391 177 397 179
rect 401 181 407 183
rect 401 179 403 181
rect 405 179 407 181
rect 401 177 407 179
rect 391 172 393 177
rect 404 172 406 177
rect 411 172 413 185
rect 435 183 437 187
rect 445 183 447 194
rect 455 191 457 194
rect 455 189 461 191
rect 455 187 457 189
rect 459 187 461 189
rect 518 205 520 209
rect 528 207 530 212
rect 538 207 540 212
rect 455 185 461 187
rect 435 181 441 183
rect 435 179 437 181
rect 439 179 441 181
rect 435 177 441 179
rect 445 181 451 183
rect 445 179 447 181
rect 449 179 451 181
rect 445 177 451 179
rect 435 172 437 177
rect 448 172 450 177
rect 455 172 457 185
rect 477 183 479 187
rect 487 183 489 194
rect 497 191 499 194
rect 497 189 503 191
rect 497 187 499 189
rect 501 187 503 189
rect 561 205 563 209
rect 571 207 573 212
rect 581 207 583 212
rect 497 185 503 187
rect 477 181 483 183
rect 477 179 479 181
rect 481 179 483 181
rect 477 177 483 179
rect 487 181 493 183
rect 487 179 489 181
rect 491 179 493 181
rect 487 177 493 179
rect 477 172 479 177
rect 490 172 492 177
rect 497 172 499 185
rect 518 183 520 187
rect 528 183 530 194
rect 538 191 540 194
rect 538 189 544 191
rect 538 187 540 189
rect 542 187 544 189
rect 601 205 603 209
rect 611 207 613 212
rect 621 207 623 212
rect 538 185 544 187
rect 518 181 524 183
rect 518 179 520 181
rect 522 179 524 181
rect 518 177 524 179
rect 528 181 534 183
rect 528 179 530 181
rect 532 179 534 181
rect 528 177 534 179
rect 518 172 520 177
rect 531 172 533 177
rect 538 172 540 185
rect 561 183 563 187
rect 571 183 573 194
rect 581 191 583 194
rect 581 189 587 191
rect 581 187 583 189
rect 585 187 587 189
rect 644 205 646 209
rect 654 207 656 212
rect 664 207 666 212
rect 581 185 587 187
rect 561 181 567 183
rect 561 179 563 181
rect 565 179 567 181
rect 561 177 567 179
rect 571 181 577 183
rect 571 179 573 181
rect 575 179 577 181
rect 571 177 577 179
rect 561 172 563 177
rect 574 172 576 177
rect 581 172 583 185
rect 601 183 603 187
rect 611 183 613 194
rect 621 191 623 194
rect 621 189 627 191
rect 621 187 623 189
rect 625 187 627 189
rect 621 185 627 187
rect 601 181 607 183
rect 601 179 603 181
rect 605 179 607 181
rect 601 177 607 179
rect 611 181 617 183
rect 611 179 613 181
rect 615 179 617 181
rect 611 177 617 179
rect 601 172 603 177
rect 614 172 616 177
rect 621 172 623 185
rect 644 183 646 187
rect 654 183 656 194
rect 664 191 666 194
rect 664 189 670 191
rect 664 187 666 189
rect 668 187 670 189
rect 664 185 670 187
rect 644 181 650 183
rect 644 179 646 181
rect 648 179 650 181
rect 644 177 650 179
rect 654 181 660 183
rect 654 179 656 181
rect 658 179 660 181
rect 654 177 660 179
rect 644 172 646 177
rect 657 172 659 177
rect 664 172 666 185
rect 49 159 51 163
rect 62 156 64 161
rect 69 156 71 161
rect 89 159 91 163
rect 102 156 104 161
rect 109 156 111 161
rect 132 159 134 163
rect 145 156 147 161
rect 152 156 154 161
rect 236 159 238 163
rect 249 156 251 161
rect 256 156 258 161
rect 278 159 280 163
rect 291 156 293 161
rect 298 156 300 161
rect 322 159 324 163
rect 335 156 337 161
rect 342 156 344 161
rect 391 159 393 163
rect 404 156 406 161
rect 411 156 413 161
rect 435 159 437 163
rect 448 156 450 161
rect 455 156 457 161
rect 477 159 479 163
rect 490 156 492 161
rect 497 156 499 161
rect 518 159 520 163
rect 531 156 533 161
rect 538 156 540 161
rect 561 159 563 163
rect 574 156 576 161
rect 581 156 583 161
rect 601 159 603 163
rect 614 156 616 161
rect 621 156 623 161
rect 644 159 646 163
rect 657 156 659 161
rect 664 156 666 161
rect -68 134 -66 138
rect -55 136 -53 141
rect -48 136 -46 141
rect 22 143 24 147
rect 33 143 35 147
rect 40 143 42 147
rect -26 134 -24 138
rect -13 136 -11 141
rect -6 136 -4 141
rect -68 120 -66 125
rect -55 120 -53 125
rect -68 118 -62 120
rect -68 116 -66 118
rect -64 116 -62 118
rect -68 114 -62 116
rect -58 118 -52 120
rect -58 116 -56 118
rect -54 116 -52 118
rect -58 114 -52 116
rect -68 110 -66 114
rect -58 103 -56 114
rect -48 112 -46 125
rect -26 120 -24 125
rect -13 120 -11 125
rect -26 118 -20 120
rect -26 116 -24 118
rect -22 116 -20 118
rect -26 114 -20 116
rect -16 118 -10 120
rect -16 116 -14 118
rect -12 116 -10 118
rect -16 114 -10 116
rect -48 110 -42 112
rect -26 110 -24 114
rect -48 108 -46 110
rect -44 108 -42 110
rect -48 106 -42 108
rect -48 103 -46 106
rect -68 88 -66 92
rect -16 103 -14 114
rect -6 112 -4 125
rect 22 120 24 129
rect 60 137 62 142
rect 70 137 72 142
rect 80 140 82 145
rect 90 143 92 147
rect 137 137 139 142
rect 156 144 178 146
rect 113 132 115 137
rect 33 120 35 123
rect 40 120 42 123
rect 60 120 62 123
rect 70 120 72 123
rect 20 118 26 120
rect 20 116 22 118
rect 24 116 26 118
rect 20 114 26 116
rect 30 118 36 120
rect 30 116 32 118
rect 34 116 36 118
rect 30 114 36 116
rect 40 118 62 120
rect 40 116 42 118
rect 44 116 49 118
rect 51 116 62 118
rect 40 114 62 116
rect 66 118 72 120
rect 66 116 68 118
rect 70 116 72 118
rect 66 114 72 116
rect 80 117 82 130
rect 90 127 92 130
rect 86 125 92 127
rect 86 123 88 125
rect 90 123 92 125
rect 149 135 151 140
rect 156 135 158 144
rect 166 135 168 140
rect 176 135 178 144
rect 203 142 205 147
rect 210 142 212 147
rect 220 145 244 147
rect 220 142 222 145
rect 86 121 92 123
rect 80 115 86 117
rect -6 110 0 112
rect 22 111 24 114
rect 32 111 34 114
rect 42 111 44 114
rect 60 111 62 114
rect 67 111 69 114
rect 80 113 82 115
rect 84 113 86 115
rect 77 111 86 113
rect -6 108 -4 110
rect -2 108 0 110
rect -6 106 0 108
rect -6 103 -4 106
rect -58 85 -56 90
rect -48 85 -46 90
rect -26 88 -24 92
rect -16 85 -14 90
rect -6 85 -4 90
rect 77 108 79 111
rect 90 108 92 121
rect 113 120 115 123
rect 137 120 139 125
rect 230 137 232 141
rect 242 140 244 145
rect 265 142 267 147
rect 272 142 274 147
rect 282 145 305 147
rect 282 142 284 145
rect 149 120 151 123
rect 156 120 158 123
rect 166 120 168 123
rect 176 120 178 123
rect 203 120 205 129
rect 210 126 212 129
rect 210 124 214 126
rect 220 124 222 129
rect 292 137 294 141
rect 242 126 244 129
rect 242 124 248 126
rect 212 120 214 124
rect 113 118 119 120
rect 113 116 115 118
rect 117 116 119 118
rect 113 114 119 116
rect 137 118 152 120
rect 137 116 139 118
rect 141 116 152 118
rect 156 117 159 120
rect 137 114 152 116
rect 113 111 115 114
rect 140 111 142 114
rect 150 111 152 114
rect 157 111 159 117
rect 163 118 169 120
rect 163 116 165 118
rect 167 116 169 118
rect 163 114 169 116
rect 176 118 183 120
rect 176 116 179 118
rect 181 116 183 118
rect 176 114 183 116
rect 202 118 208 120
rect 202 116 204 118
rect 206 116 208 118
rect 202 114 208 116
rect 212 118 218 120
rect 212 116 214 118
rect 216 116 218 118
rect 230 116 232 124
rect 242 122 244 124
rect 246 122 248 124
rect 242 120 248 122
rect 265 120 267 129
rect 272 120 274 129
rect 282 124 284 129
rect 303 134 305 145
rect 355 137 357 142
rect 374 144 396 146
rect 292 121 294 124
rect 331 132 333 137
rect 367 135 369 140
rect 374 135 376 144
rect 384 135 386 140
rect 394 135 396 144
rect 421 142 423 147
rect 428 142 430 147
rect 438 145 462 147
rect 438 142 440 145
rect 252 118 258 120
rect 252 116 254 118
rect 256 116 258 118
rect 212 114 218 116
rect 222 114 258 116
rect 262 118 268 120
rect 262 116 264 118
rect 266 116 268 118
rect 262 114 268 116
rect 272 118 278 120
rect 272 116 274 118
rect 276 116 278 118
rect 290 119 296 121
rect 290 117 292 119
rect 294 117 296 119
rect 272 114 278 116
rect 282 115 296 117
rect 167 111 169 114
rect 177 111 179 114
rect 202 111 204 114
rect 212 111 214 114
rect 222 111 224 114
rect 262 111 264 114
rect 272 111 274 114
rect 282 111 284 115
rect 77 90 79 95
rect 22 79 24 83
rect 32 79 34 83
rect 42 79 44 83
rect 60 81 62 86
rect 67 81 69 86
rect 113 88 115 93
rect 90 79 92 83
rect 140 79 142 84
rect 150 79 152 84
rect 157 79 159 84
rect 167 79 169 84
rect 177 79 179 84
rect 238 104 244 106
rect 238 102 240 104
rect 242 102 244 104
rect 232 100 244 102
rect 232 97 234 100
rect 242 97 244 100
rect 303 109 305 123
rect 331 120 333 123
rect 355 120 357 125
rect 448 137 450 141
rect 460 140 462 145
rect 483 142 485 147
rect 490 142 492 147
rect 500 145 523 147
rect 500 142 502 145
rect 367 120 369 123
rect 374 120 376 123
rect 384 120 386 123
rect 394 120 396 123
rect 421 120 423 129
rect 428 126 430 129
rect 428 124 432 126
rect 438 124 440 129
rect 510 137 512 141
rect 460 126 462 129
rect 460 124 466 126
rect 430 120 432 124
rect 331 118 337 120
rect 331 116 333 118
rect 335 116 337 118
rect 331 114 337 116
rect 355 118 370 120
rect 355 116 357 118
rect 359 116 370 118
rect 374 117 377 120
rect 355 114 370 116
rect 313 111 319 113
rect 331 111 333 114
rect 358 111 360 114
rect 368 111 370 114
rect 375 111 377 117
rect 381 118 387 120
rect 381 116 383 118
rect 385 116 387 118
rect 381 114 387 116
rect 394 118 401 120
rect 394 116 397 118
rect 399 116 401 118
rect 394 114 401 116
rect 420 118 426 120
rect 420 116 422 118
rect 424 116 426 118
rect 420 114 426 116
rect 430 118 436 120
rect 430 116 432 118
rect 434 116 436 118
rect 448 116 450 124
rect 460 122 462 124
rect 464 122 466 124
rect 460 120 466 122
rect 483 120 485 129
rect 490 120 492 129
rect 500 124 502 129
rect 521 134 523 145
rect 560 143 562 147
rect 571 143 573 147
rect 578 143 580 147
rect 510 121 512 124
rect 470 118 476 120
rect 470 116 472 118
rect 474 116 476 118
rect 430 114 436 116
rect 440 114 476 116
rect 480 118 486 120
rect 480 116 482 118
rect 484 116 486 118
rect 480 114 486 116
rect 490 118 496 120
rect 490 116 492 118
rect 494 116 496 118
rect 508 119 514 121
rect 508 117 510 119
rect 512 117 514 119
rect 490 114 496 116
rect 500 115 514 117
rect 385 111 387 114
rect 395 111 397 114
rect 420 111 422 114
rect 430 111 432 114
rect 440 111 442 114
rect 480 111 482 114
rect 490 111 492 114
rect 500 111 502 115
rect 313 109 315 111
rect 317 109 319 111
rect 293 107 319 109
rect 293 104 295 107
rect 303 104 305 107
rect 293 86 295 90
rect 303 86 305 90
rect 331 88 333 93
rect 202 79 204 83
rect 212 79 214 83
rect 222 79 224 83
rect 232 79 234 83
rect 242 79 244 83
rect 262 79 264 83
rect 272 79 274 83
rect 282 79 284 83
rect 358 79 360 84
rect 368 79 370 84
rect 375 79 377 84
rect 385 79 387 84
rect 395 79 397 84
rect 456 104 462 106
rect 456 102 458 104
rect 460 102 462 104
rect 450 100 462 102
rect 450 97 452 100
rect 460 97 462 100
rect 521 109 523 123
rect 560 120 562 129
rect 598 137 600 142
rect 608 137 610 142
rect 618 140 620 145
rect 628 143 630 147
rect 571 120 573 123
rect 578 120 580 123
rect 598 120 600 123
rect 608 120 610 123
rect 558 118 564 120
rect 558 116 560 118
rect 562 116 564 118
rect 558 114 564 116
rect 568 118 574 120
rect 568 116 570 118
rect 572 116 574 118
rect 568 114 574 116
rect 578 118 600 120
rect 578 116 580 118
rect 582 116 587 118
rect 589 116 600 118
rect 578 114 600 116
rect 604 118 610 120
rect 604 116 606 118
rect 608 116 610 118
rect 604 114 610 116
rect 618 117 620 130
rect 628 127 630 130
rect 624 125 630 127
rect 624 123 626 125
rect 628 123 630 125
rect 624 121 630 123
rect 618 115 624 117
rect 531 111 537 113
rect 560 111 562 114
rect 570 111 572 114
rect 580 111 582 114
rect 598 111 600 114
rect 605 111 607 114
rect 618 113 620 115
rect 622 113 624 115
rect 615 111 624 113
rect 531 109 533 111
rect 535 109 537 111
rect 511 107 537 109
rect 511 104 513 107
rect 521 104 523 107
rect 511 86 513 90
rect 521 86 523 90
rect 420 79 422 83
rect 430 79 432 83
rect 440 79 442 83
rect 450 79 452 83
rect 460 79 462 83
rect 480 79 482 83
rect 490 79 492 83
rect 500 79 502 83
rect 615 108 617 111
rect 628 108 630 121
rect 615 90 617 95
rect 560 79 562 83
rect 570 79 572 83
rect 580 79 582 83
rect 598 81 600 86
rect 605 81 607 86
rect 628 79 630 83
rect -114 70 -112 75
rect -104 70 -102 75
rect -97 70 -95 75
rect -87 70 -85 75
rect -77 70 -75 75
rect -52 71 -50 75
rect -42 71 -40 75
rect -32 71 -30 75
rect -22 71 -20 75
rect -12 71 -10 75
rect 8 71 10 75
rect 18 71 20 75
rect 28 71 30 75
rect -185 62 -183 66
rect -175 64 -173 69
rect -165 64 -163 69
rect -141 61 -139 66
rect -185 40 -183 44
rect -175 40 -173 51
rect -165 48 -163 51
rect -165 46 -159 48
rect -165 44 -163 46
rect -161 44 -159 46
rect -165 42 -159 44
rect -22 54 -20 57
rect -12 54 -10 57
rect -22 52 -10 54
rect -16 50 -14 52
rect -12 50 -10 52
rect -16 48 -10 50
rect 104 70 106 75
rect 114 70 116 75
rect 121 70 123 75
rect 131 70 133 75
rect 141 70 143 75
rect 166 71 168 75
rect 176 71 178 75
rect 186 71 188 75
rect 196 71 198 75
rect 206 71 208 75
rect 226 71 228 75
rect 236 71 238 75
rect 246 71 248 75
rect 39 64 41 68
rect 49 64 51 68
rect 77 61 79 66
rect 39 47 41 50
rect 49 47 51 50
rect 39 45 65 47
rect -185 38 -179 40
rect -185 36 -183 38
rect -181 36 -179 38
rect -185 34 -179 36
rect -175 38 -169 40
rect -175 36 -173 38
rect -171 36 -169 38
rect -175 34 -169 36
rect -185 29 -183 34
rect -172 29 -170 34
rect -165 29 -163 42
rect -141 40 -139 43
rect -114 40 -112 43
rect -104 40 -102 43
rect -141 38 -135 40
rect -141 36 -139 38
rect -137 36 -135 38
rect -141 34 -135 36
rect -117 38 -102 40
rect -117 36 -115 38
rect -113 36 -102 38
rect -97 37 -95 43
rect -87 40 -85 43
rect -77 40 -75 43
rect -52 40 -50 43
rect -42 40 -40 43
rect -32 40 -30 43
rect 8 40 10 43
rect 18 40 20 43
rect -117 34 -102 36
rect -98 34 -95 37
rect -91 38 -85 40
rect -91 36 -89 38
rect -87 36 -85 38
rect -91 34 -85 36
rect -78 38 -71 40
rect -78 36 -75 38
rect -73 36 -71 38
rect -78 34 -71 36
rect -52 38 -46 40
rect -52 36 -50 38
rect -48 36 -46 38
rect -52 34 -46 36
rect -42 38 -36 40
rect -32 38 4 40
rect -42 36 -40 38
rect -38 36 -36 38
rect -42 34 -36 36
rect -141 31 -139 34
rect -185 16 -183 20
rect -117 29 -115 34
rect -105 31 -103 34
rect -98 31 -96 34
rect -88 31 -86 34
rect -78 31 -76 34
rect -172 13 -170 18
rect -165 13 -163 18
rect -141 17 -139 22
rect -51 25 -49 34
rect -42 30 -40 34
rect -24 30 -22 38
rect -2 36 0 38
rect 2 36 4 38
rect -2 34 4 36
rect 8 38 14 40
rect 8 36 10 38
rect 12 36 14 38
rect 8 34 14 36
rect 18 38 24 40
rect 18 36 20 38
rect 22 36 24 38
rect 28 39 30 43
rect 28 37 42 39
rect 18 34 24 36
rect 36 35 38 37
rect 40 35 42 37
rect -12 32 -6 34
rect -12 30 -10 32
rect -8 30 -6 32
rect -44 28 -40 30
rect -44 25 -42 28
rect -34 25 -32 30
rect -117 12 -115 17
rect -105 14 -103 19
rect -98 10 -96 19
rect -88 14 -86 19
rect -78 10 -76 19
rect -98 8 -76 10
rect -12 28 -6 30
rect -12 25 -10 28
rect 11 25 13 34
rect 18 25 20 34
rect 36 33 42 35
rect 38 30 40 33
rect 49 31 51 45
rect 59 43 61 45
rect 63 43 65 45
rect 196 54 198 57
rect 206 54 208 57
rect 196 52 208 54
rect 202 50 204 52
rect 206 50 208 52
rect 202 48 208 50
rect 324 70 326 75
rect 334 70 336 75
rect 341 70 343 75
rect 351 70 353 75
rect 361 70 363 75
rect 386 71 388 75
rect 396 71 398 75
rect 406 71 408 75
rect 416 71 418 75
rect 426 71 428 75
rect 446 71 448 75
rect 456 71 458 75
rect 466 71 468 75
rect 257 64 259 68
rect 267 64 269 68
rect 297 61 299 66
rect 257 47 259 50
rect 267 47 269 50
rect 257 45 283 47
rect 59 41 65 43
rect 77 40 79 43
rect 104 40 106 43
rect 114 40 116 43
rect 77 38 83 40
rect 77 36 79 38
rect 81 36 83 38
rect 77 34 83 36
rect 101 38 116 40
rect 101 36 103 38
rect 105 36 116 38
rect 121 37 123 43
rect 131 40 133 43
rect 141 40 143 43
rect 166 40 168 43
rect 176 40 178 43
rect 186 40 188 43
rect 226 40 228 43
rect 236 40 238 43
rect 101 34 116 36
rect 120 34 123 37
rect 127 38 133 40
rect 127 36 129 38
rect 131 36 133 38
rect 127 34 133 36
rect 140 38 147 40
rect 140 36 143 38
rect 145 36 147 38
rect 140 34 147 36
rect 166 38 172 40
rect 166 36 168 38
rect 170 36 172 38
rect 166 34 172 36
rect 176 38 182 40
rect 186 38 222 40
rect 176 36 178 38
rect 180 36 182 38
rect 176 34 182 36
rect 77 31 79 34
rect 28 25 30 30
rect -24 13 -22 17
rect -51 7 -49 12
rect -44 7 -42 12
rect -34 9 -32 12
rect -12 9 -10 14
rect -34 7 -10 9
rect 101 29 103 34
rect 113 31 115 34
rect 120 31 122 34
rect 130 31 132 34
rect 140 31 142 34
rect 38 13 40 17
rect 11 7 13 12
rect 18 7 20 12
rect 28 9 30 12
rect 49 9 51 20
rect 77 17 79 22
rect 167 25 169 34
rect 176 30 178 34
rect 194 30 196 38
rect 216 36 218 38
rect 220 36 222 38
rect 216 34 222 36
rect 226 38 232 40
rect 226 36 228 38
rect 230 36 232 38
rect 226 34 232 36
rect 236 38 242 40
rect 236 36 238 38
rect 240 36 242 38
rect 246 39 248 43
rect 246 37 260 39
rect 236 34 242 36
rect 254 35 256 37
rect 258 35 260 37
rect 206 32 212 34
rect 206 30 208 32
rect 210 30 212 32
rect 174 28 178 30
rect 174 25 176 28
rect 184 25 186 30
rect 28 7 51 9
rect 101 12 103 17
rect 113 14 115 19
rect 120 10 122 19
rect 130 14 132 19
rect 140 10 142 19
rect 120 8 142 10
rect 206 28 212 30
rect 206 25 208 28
rect 229 25 231 34
rect 236 25 238 34
rect 254 33 260 35
rect 256 30 258 33
rect 267 31 269 45
rect 277 43 279 45
rect 281 43 283 45
rect 416 54 418 57
rect 426 54 428 57
rect 416 52 428 54
rect 422 50 424 52
rect 426 50 428 52
rect 422 48 428 50
rect 519 71 521 75
rect 529 71 531 75
rect 539 71 541 75
rect 477 64 479 68
rect 487 64 489 68
rect 477 47 479 50
rect 487 47 489 50
rect 477 45 503 47
rect 277 41 283 43
rect 297 40 299 43
rect 324 40 326 43
rect 334 40 336 43
rect 297 38 303 40
rect 297 36 299 38
rect 301 36 303 38
rect 297 34 303 36
rect 321 38 336 40
rect 321 36 323 38
rect 325 36 336 38
rect 341 37 343 43
rect 351 40 353 43
rect 361 40 363 43
rect 386 40 388 43
rect 396 40 398 43
rect 406 40 408 43
rect 446 40 448 43
rect 456 40 458 43
rect 321 34 336 36
rect 340 34 343 37
rect 347 38 353 40
rect 347 36 349 38
rect 351 36 353 38
rect 347 34 353 36
rect 360 38 367 40
rect 360 36 363 38
rect 365 36 367 38
rect 360 34 367 36
rect 386 38 392 40
rect 386 36 388 38
rect 390 36 392 38
rect 386 34 392 36
rect 396 38 402 40
rect 406 38 442 40
rect 396 36 398 38
rect 400 36 402 38
rect 396 34 402 36
rect 297 31 299 34
rect 246 25 248 30
rect 194 13 196 17
rect 167 7 169 12
rect 174 7 176 12
rect 184 9 186 12
rect 206 9 208 14
rect 184 7 208 9
rect 321 29 323 34
rect 333 31 335 34
rect 340 31 342 34
rect 350 31 352 34
rect 360 31 362 34
rect 256 13 258 17
rect 229 7 231 12
rect 236 7 238 12
rect 246 9 248 12
rect 267 9 269 20
rect 297 17 299 22
rect 387 25 389 34
rect 396 30 398 34
rect 414 30 416 38
rect 436 36 438 38
rect 440 36 442 38
rect 436 34 442 36
rect 446 38 452 40
rect 446 36 448 38
rect 450 36 452 38
rect 446 34 452 36
rect 456 38 462 40
rect 456 36 458 38
rect 460 36 462 38
rect 466 39 468 43
rect 466 37 480 39
rect 456 34 462 36
rect 474 35 476 37
rect 478 35 480 37
rect 426 32 432 34
rect 426 30 428 32
rect 430 30 432 32
rect 394 28 398 30
rect 394 25 396 28
rect 404 25 406 30
rect 246 7 269 9
rect 321 12 323 17
rect 333 14 335 19
rect 340 10 342 19
rect 350 14 352 19
rect 360 10 362 19
rect 340 8 362 10
rect 426 28 432 30
rect 426 25 428 28
rect 449 25 451 34
rect 456 25 458 34
rect 474 33 480 35
rect 476 30 478 33
rect 487 31 489 45
rect 497 43 499 45
rect 501 43 503 45
rect 557 68 559 73
rect 564 68 566 73
rect 587 71 589 75
rect 574 59 576 64
rect 574 43 576 46
rect 497 41 503 43
rect 519 40 521 43
rect 529 40 531 43
rect 539 40 541 43
rect 557 40 559 43
rect 564 40 566 43
rect 574 41 583 43
rect 517 38 523 40
rect 517 36 519 38
rect 521 36 523 38
rect 517 34 523 36
rect 527 38 533 40
rect 527 36 529 38
rect 531 36 533 38
rect 527 34 533 36
rect 537 38 559 40
rect 537 36 539 38
rect 541 36 546 38
rect 548 36 559 38
rect 537 34 559 36
rect 563 38 569 40
rect 563 36 565 38
rect 567 36 569 38
rect 563 34 569 36
rect 466 25 468 30
rect 414 13 416 17
rect 387 7 389 12
rect 394 7 396 12
rect 404 9 406 12
rect 426 9 428 14
rect 404 7 428 9
rect 519 25 521 34
rect 530 31 532 34
rect 537 31 539 34
rect 557 31 559 34
rect 567 31 569 34
rect 577 39 579 41
rect 581 39 583 41
rect 577 37 583 39
rect 476 13 478 17
rect 449 7 451 12
rect 456 7 458 12
rect 466 9 468 12
rect 487 9 489 20
rect 466 7 489 9
rect 577 24 579 37
rect 587 33 589 46
rect 583 31 589 33
rect 583 29 585 31
rect 587 29 589 31
rect 583 27 589 29
rect 587 24 589 27
rect 557 12 559 17
rect 567 12 569 17
rect 519 7 521 11
rect 530 7 532 11
rect 537 7 539 11
rect 577 9 579 14
rect 587 7 589 11
rect -179 -7 -177 -2
rect -160 0 -138 2
rect -203 -12 -201 -7
rect -167 -9 -165 -4
rect -160 -9 -158 0
rect -150 -9 -148 -4
rect -140 -9 -138 0
rect -113 -2 -111 3
rect -106 -2 -104 3
rect -96 1 -72 3
rect -96 -2 -94 1
rect -203 -24 -201 -21
rect -179 -24 -177 -19
rect -86 -7 -84 -3
rect -74 -4 -72 1
rect -51 -2 -49 3
rect -44 -2 -42 3
rect -34 1 -11 3
rect -34 -2 -32 1
rect -167 -24 -165 -21
rect -160 -24 -158 -21
rect -150 -24 -148 -21
rect -140 -24 -138 -21
rect -113 -24 -111 -15
rect -106 -18 -104 -15
rect -106 -20 -102 -18
rect -96 -20 -94 -15
rect -24 -7 -22 -3
rect -74 -18 -72 -15
rect -74 -20 -68 -18
rect -104 -24 -102 -20
rect -203 -26 -197 -24
rect -203 -28 -201 -26
rect -199 -28 -197 -26
rect -203 -30 -197 -28
rect -179 -26 -164 -24
rect -179 -28 -177 -26
rect -175 -28 -164 -26
rect -160 -27 -157 -24
rect -179 -30 -164 -28
rect -203 -33 -201 -30
rect -176 -33 -174 -30
rect -166 -33 -164 -30
rect -159 -33 -157 -27
rect -153 -26 -147 -24
rect -153 -28 -151 -26
rect -149 -28 -147 -26
rect -153 -30 -147 -28
rect -140 -26 -133 -24
rect -140 -28 -137 -26
rect -135 -28 -133 -26
rect -140 -30 -133 -28
rect -114 -26 -108 -24
rect -114 -28 -112 -26
rect -110 -28 -108 -26
rect -114 -30 -108 -28
rect -104 -26 -98 -24
rect -104 -28 -102 -26
rect -100 -28 -98 -26
rect -86 -28 -84 -20
rect -74 -22 -72 -20
rect -70 -22 -68 -20
rect -74 -24 -68 -22
rect -51 -24 -49 -15
rect -44 -24 -42 -15
rect -34 -20 -32 -15
rect -13 -10 -11 1
rect 41 -7 43 -2
rect 60 0 82 2
rect -24 -23 -22 -20
rect 17 -12 19 -7
rect 53 -9 55 -4
rect 60 -9 62 0
rect 70 -9 72 -4
rect 80 -9 82 0
rect 107 -2 109 3
rect 114 -2 116 3
rect 124 1 148 3
rect 124 -2 126 1
rect -64 -26 -58 -24
rect -64 -28 -62 -26
rect -60 -28 -58 -26
rect -104 -30 -98 -28
rect -94 -30 -58 -28
rect -54 -26 -48 -24
rect -54 -28 -52 -26
rect -50 -28 -48 -26
rect -54 -30 -48 -28
rect -44 -26 -38 -24
rect -44 -28 -42 -26
rect -40 -28 -38 -26
rect -26 -25 -20 -23
rect -26 -27 -24 -25
rect -22 -27 -20 -25
rect -44 -30 -38 -28
rect -34 -29 -20 -27
rect -149 -33 -147 -30
rect -139 -33 -137 -30
rect -114 -33 -112 -30
rect -104 -33 -102 -30
rect -94 -33 -92 -30
rect -54 -33 -52 -30
rect -44 -33 -42 -30
rect -34 -33 -32 -29
rect -203 -56 -201 -51
rect -176 -65 -174 -60
rect -166 -65 -164 -60
rect -159 -65 -157 -60
rect -149 -65 -147 -60
rect -139 -65 -137 -60
rect -78 -40 -72 -38
rect -78 -42 -76 -40
rect -74 -42 -72 -40
rect -84 -44 -72 -42
rect -84 -47 -82 -44
rect -74 -47 -72 -44
rect -13 -35 -11 -21
rect 17 -24 19 -21
rect 41 -24 43 -19
rect 134 -7 136 -3
rect 146 -4 148 1
rect 169 -2 171 3
rect 176 -2 178 3
rect 186 1 209 3
rect 186 -2 188 1
rect 53 -24 55 -21
rect 60 -24 62 -21
rect 70 -24 72 -21
rect 80 -24 82 -21
rect 107 -24 109 -15
rect 114 -18 116 -15
rect 114 -20 118 -18
rect 124 -20 126 -15
rect 196 -7 198 -3
rect 146 -18 148 -15
rect 146 -20 152 -18
rect 116 -24 118 -20
rect 17 -26 23 -24
rect 17 -28 19 -26
rect 21 -28 23 -26
rect 17 -30 23 -28
rect 41 -26 56 -24
rect 41 -28 43 -26
rect 45 -28 56 -26
rect 60 -27 63 -24
rect 41 -30 56 -28
rect -3 -33 3 -31
rect 17 -33 19 -30
rect 44 -33 46 -30
rect 54 -33 56 -30
rect 61 -33 63 -27
rect 67 -26 73 -24
rect 67 -28 69 -26
rect 71 -28 73 -26
rect 67 -30 73 -28
rect 80 -26 87 -24
rect 80 -28 83 -26
rect 85 -28 87 -26
rect 80 -30 87 -28
rect 106 -26 112 -24
rect 106 -28 108 -26
rect 110 -28 112 -26
rect 106 -30 112 -28
rect 116 -26 122 -24
rect 116 -28 118 -26
rect 120 -28 122 -26
rect 134 -28 136 -20
rect 146 -22 148 -20
rect 150 -22 152 -20
rect 146 -24 152 -22
rect 169 -24 171 -15
rect 176 -24 178 -15
rect 186 -20 188 -15
rect 207 -10 209 1
rect 258 -7 260 -2
rect 277 0 299 2
rect 196 -23 198 -20
rect 234 -12 236 -7
rect 270 -9 272 -4
rect 277 -9 279 0
rect 287 -9 289 -4
rect 297 -9 299 0
rect 324 -2 326 3
rect 331 -2 333 3
rect 341 1 365 3
rect 341 -2 343 1
rect 156 -26 162 -24
rect 156 -28 158 -26
rect 160 -28 162 -26
rect 116 -30 122 -28
rect 126 -30 162 -28
rect 166 -26 172 -24
rect 166 -28 168 -26
rect 170 -28 172 -26
rect 166 -30 172 -28
rect 176 -26 182 -24
rect 176 -28 178 -26
rect 180 -28 182 -26
rect 194 -25 200 -23
rect 194 -27 196 -25
rect 198 -27 200 -25
rect 176 -30 182 -28
rect 186 -29 200 -27
rect 71 -33 73 -30
rect 81 -33 83 -30
rect 106 -33 108 -30
rect 116 -33 118 -30
rect 126 -33 128 -30
rect 166 -33 168 -30
rect 176 -33 178 -30
rect 186 -33 188 -29
rect -3 -35 -1 -33
rect 1 -35 3 -33
rect -23 -37 3 -35
rect -23 -40 -21 -37
rect -13 -40 -11 -37
rect -23 -58 -21 -54
rect -13 -58 -11 -54
rect 17 -56 19 -51
rect -114 -65 -112 -61
rect -104 -65 -102 -61
rect -94 -65 -92 -61
rect -84 -65 -82 -61
rect -74 -65 -72 -61
rect -54 -65 -52 -61
rect -44 -65 -42 -61
rect -34 -65 -32 -61
rect 44 -65 46 -60
rect 54 -65 56 -60
rect 61 -65 63 -60
rect 71 -65 73 -60
rect 81 -65 83 -60
rect 142 -40 148 -38
rect 142 -42 144 -40
rect 146 -42 148 -40
rect 136 -44 148 -42
rect 136 -47 138 -44
rect 146 -47 148 -44
rect 207 -35 209 -21
rect 234 -24 236 -21
rect 258 -24 260 -19
rect 351 -7 353 -3
rect 363 -4 365 1
rect 386 -2 388 3
rect 393 -2 395 3
rect 403 1 426 3
rect 403 -2 405 1
rect 270 -24 272 -21
rect 277 -24 279 -21
rect 287 -24 289 -21
rect 297 -24 299 -21
rect 324 -24 326 -15
rect 331 -18 333 -15
rect 331 -20 335 -18
rect 341 -20 343 -15
rect 413 -7 415 -3
rect 363 -18 365 -15
rect 363 -20 369 -18
rect 333 -24 335 -20
rect 234 -26 240 -24
rect 234 -28 236 -26
rect 238 -28 240 -26
rect 234 -30 240 -28
rect 258 -26 273 -24
rect 258 -28 260 -26
rect 262 -28 273 -26
rect 277 -27 280 -24
rect 258 -30 273 -28
rect 217 -33 223 -31
rect 234 -33 236 -30
rect 261 -33 263 -30
rect 271 -33 273 -30
rect 278 -33 280 -27
rect 284 -26 290 -24
rect 284 -28 286 -26
rect 288 -28 290 -26
rect 284 -30 290 -28
rect 297 -26 304 -24
rect 297 -28 300 -26
rect 302 -28 304 -26
rect 297 -30 304 -28
rect 323 -26 329 -24
rect 323 -28 325 -26
rect 327 -28 329 -26
rect 323 -30 329 -28
rect 333 -26 339 -24
rect 333 -28 335 -26
rect 337 -28 339 -26
rect 351 -28 353 -20
rect 363 -22 365 -20
rect 367 -22 369 -20
rect 363 -24 369 -22
rect 386 -24 388 -15
rect 393 -24 395 -15
rect 403 -20 405 -15
rect 424 -10 426 1
rect 462 -1 464 3
rect 473 -1 475 3
rect 480 -1 482 3
rect 413 -23 415 -20
rect 373 -26 379 -24
rect 373 -28 375 -26
rect 377 -28 379 -26
rect 333 -30 339 -28
rect 343 -30 379 -28
rect 383 -26 389 -24
rect 383 -28 385 -26
rect 387 -28 389 -26
rect 383 -30 389 -28
rect 393 -26 399 -24
rect 393 -28 395 -26
rect 397 -28 399 -26
rect 411 -25 417 -23
rect 411 -27 413 -25
rect 415 -27 417 -25
rect 393 -30 399 -28
rect 403 -29 417 -27
rect 288 -33 290 -30
rect 298 -33 300 -30
rect 323 -33 325 -30
rect 333 -33 335 -30
rect 343 -33 345 -30
rect 383 -33 385 -30
rect 393 -33 395 -30
rect 403 -33 405 -29
rect 217 -35 219 -33
rect 221 -35 223 -33
rect 197 -37 223 -35
rect 197 -40 199 -37
rect 207 -40 209 -37
rect 197 -58 199 -54
rect 207 -58 209 -54
rect 234 -56 236 -51
rect 106 -65 108 -61
rect 116 -65 118 -61
rect 126 -65 128 -61
rect 136 -65 138 -61
rect 146 -65 148 -61
rect 166 -65 168 -61
rect 176 -65 178 -61
rect 186 -65 188 -61
rect 261 -65 263 -60
rect 271 -65 273 -60
rect 278 -65 280 -60
rect 288 -65 290 -60
rect 298 -65 300 -60
rect 359 -40 365 -38
rect 359 -42 361 -40
rect 363 -42 365 -40
rect 353 -44 365 -42
rect 353 -47 355 -44
rect 363 -47 365 -44
rect 424 -35 426 -21
rect 462 -24 464 -15
rect 500 -7 502 -2
rect 510 -7 512 -2
rect 520 -4 522 1
rect 530 -1 532 3
rect 473 -24 475 -21
rect 480 -24 482 -21
rect 500 -24 502 -21
rect 510 -24 512 -21
rect 460 -26 466 -24
rect 460 -28 462 -26
rect 464 -28 466 -26
rect 460 -30 466 -28
rect 470 -26 476 -24
rect 470 -28 472 -26
rect 474 -28 476 -26
rect 470 -30 476 -28
rect 480 -26 502 -24
rect 480 -28 482 -26
rect 484 -28 489 -26
rect 491 -28 502 -26
rect 480 -30 502 -28
rect 506 -26 512 -24
rect 506 -28 508 -26
rect 510 -28 512 -26
rect 506 -30 512 -28
rect 520 -27 522 -14
rect 530 -17 532 -14
rect 526 -19 532 -17
rect 526 -21 528 -19
rect 530 -21 532 -19
rect 526 -23 532 -21
rect 520 -29 526 -27
rect 434 -33 440 -31
rect 462 -33 464 -30
rect 472 -33 474 -30
rect 482 -33 484 -30
rect 500 -33 502 -30
rect 507 -33 509 -30
rect 520 -31 522 -29
rect 524 -31 526 -29
rect 517 -33 526 -31
rect 434 -35 436 -33
rect 438 -35 440 -33
rect 414 -37 440 -35
rect 414 -40 416 -37
rect 424 -40 426 -37
rect 414 -58 416 -54
rect 424 -58 426 -54
rect 323 -65 325 -61
rect 333 -65 335 -61
rect 343 -65 345 -61
rect 353 -65 355 -61
rect 363 -65 365 -61
rect 383 -65 385 -61
rect 393 -65 395 -61
rect 403 -65 405 -61
rect 517 -36 519 -33
rect 530 -36 532 -23
rect 517 -54 519 -49
rect 462 -65 464 -61
rect 472 -65 474 -61
rect 482 -65 484 -61
rect 500 -63 502 -58
rect 507 -63 509 -58
rect 530 -65 532 -61
<< ndif >>
rect 44 169 49 172
rect 42 167 49 169
rect 42 165 44 167
rect 46 165 49 167
rect 42 163 49 165
rect 51 163 62 172
rect 53 161 62 163
rect 64 161 69 172
rect 71 167 76 172
rect 84 169 89 172
rect 82 167 89 169
rect 71 165 78 167
rect 71 163 74 165
rect 76 163 78 165
rect 82 165 84 167
rect 86 165 89 167
rect 82 163 89 165
rect 91 163 102 172
rect 71 161 78 163
rect 53 155 60 161
rect 93 161 102 163
rect 104 161 109 172
rect 111 167 116 172
rect 127 169 132 172
rect 125 167 132 169
rect 111 165 118 167
rect 111 163 114 165
rect 116 163 118 165
rect 125 165 127 167
rect 129 165 132 167
rect 125 163 132 165
rect 134 163 145 172
rect 111 161 118 163
rect 53 153 55 155
rect 57 153 60 155
rect 53 151 60 153
rect 93 155 100 161
rect 136 161 145 163
rect 147 161 152 172
rect 154 167 159 172
rect 231 169 236 172
rect 229 167 236 169
rect 154 165 161 167
rect 154 163 157 165
rect 159 163 161 165
rect 229 165 231 167
rect 233 165 236 167
rect 229 163 236 165
rect 238 163 249 172
rect 154 161 161 163
rect 93 153 95 155
rect 97 153 100 155
rect 93 151 100 153
rect 136 155 143 161
rect 240 161 249 163
rect 251 161 256 172
rect 258 167 263 172
rect 273 169 278 172
rect 271 167 278 169
rect 258 165 265 167
rect 258 163 261 165
rect 263 163 265 165
rect 271 165 273 167
rect 275 165 278 167
rect 271 163 278 165
rect 280 163 291 172
rect 258 161 265 163
rect 136 153 138 155
rect 140 153 143 155
rect 136 151 143 153
rect 240 155 247 161
rect 282 161 291 163
rect 293 161 298 172
rect 300 167 305 172
rect 317 169 322 172
rect 315 167 322 169
rect 300 165 307 167
rect 300 163 303 165
rect 305 163 307 165
rect 315 165 317 167
rect 319 165 322 167
rect 315 163 322 165
rect 324 163 335 172
rect 300 161 307 163
rect 240 153 242 155
rect 244 153 247 155
rect 240 151 247 153
rect 282 155 289 161
rect 326 161 335 163
rect 337 161 342 172
rect 344 167 349 172
rect 386 169 391 172
rect 384 167 391 169
rect 344 165 351 167
rect 344 163 347 165
rect 349 163 351 165
rect 384 165 386 167
rect 388 165 391 167
rect 384 163 391 165
rect 393 163 404 172
rect 344 161 351 163
rect 282 153 284 155
rect 286 153 289 155
rect 282 151 289 153
rect 326 155 333 161
rect 395 161 404 163
rect 406 161 411 172
rect 413 167 418 172
rect 430 169 435 172
rect 428 167 435 169
rect 413 165 420 167
rect 413 163 416 165
rect 418 163 420 165
rect 428 165 430 167
rect 432 165 435 167
rect 428 163 435 165
rect 437 163 448 172
rect 413 161 420 163
rect 326 153 328 155
rect 330 153 333 155
rect 326 151 333 153
rect 395 155 402 161
rect 439 161 448 163
rect 450 161 455 172
rect 457 167 462 172
rect 472 169 477 172
rect 470 167 477 169
rect 457 165 464 167
rect 457 163 460 165
rect 462 163 464 165
rect 470 165 472 167
rect 474 165 477 167
rect 470 163 477 165
rect 479 163 490 172
rect 457 161 464 163
rect 395 153 397 155
rect 399 153 402 155
rect 395 151 402 153
rect 439 155 446 161
rect 481 161 490 163
rect 492 161 497 172
rect 499 167 504 172
rect 513 169 518 172
rect 511 167 518 169
rect 499 165 506 167
rect 499 163 502 165
rect 504 163 506 165
rect 511 165 513 167
rect 515 165 518 167
rect 511 163 518 165
rect 520 163 531 172
rect 499 161 506 163
rect 439 153 441 155
rect 443 153 446 155
rect 439 151 446 153
rect 481 155 488 161
rect 522 161 531 163
rect 533 161 538 172
rect 540 167 545 172
rect 556 169 561 172
rect 554 167 561 169
rect 540 165 547 167
rect 540 163 543 165
rect 545 163 547 165
rect 554 165 556 167
rect 558 165 561 167
rect 554 163 561 165
rect 563 163 574 172
rect 540 161 547 163
rect 481 153 483 155
rect 485 153 488 155
rect 481 151 488 153
rect 522 155 529 161
rect 565 161 574 163
rect 576 161 581 172
rect 583 167 588 172
rect 596 169 601 172
rect 594 167 601 169
rect 583 165 590 167
rect 583 163 586 165
rect 588 163 590 165
rect 594 165 596 167
rect 598 165 601 167
rect 594 163 601 165
rect 603 163 614 172
rect 583 161 590 163
rect 522 153 524 155
rect 526 153 529 155
rect 522 151 529 153
rect 565 155 572 161
rect 605 161 614 163
rect 616 161 621 172
rect 623 167 628 172
rect 639 169 644 172
rect 637 167 644 169
rect 623 165 630 167
rect 623 163 626 165
rect 628 163 630 165
rect 637 165 639 167
rect 641 165 644 167
rect 637 163 644 165
rect 646 163 657 172
rect 623 161 630 163
rect 565 153 567 155
rect 569 153 572 155
rect 565 151 572 153
rect 605 155 612 161
rect 648 161 657 163
rect 659 161 664 172
rect 666 167 671 172
rect 666 165 673 167
rect 666 163 669 165
rect 671 163 673 165
rect 666 161 673 163
rect 605 153 607 155
rect 609 153 612 155
rect 605 151 612 153
rect 648 155 655 161
rect 648 153 650 155
rect 652 153 655 155
rect 648 151 655 153
rect -64 144 -57 146
rect -64 142 -62 144
rect -60 142 -57 144
rect -64 136 -57 142
rect -22 144 -15 146
rect -22 142 -20 144
rect -18 142 -15 144
rect -64 134 -55 136
rect -75 132 -68 134
rect -75 130 -73 132
rect -71 130 -68 132
rect -75 128 -68 130
rect -73 125 -68 128
rect -66 125 -55 134
rect -53 125 -48 136
rect -46 134 -39 136
rect -22 136 -15 142
rect 17 136 22 143
rect -22 134 -13 136
rect -46 132 -43 134
rect -41 132 -39 134
rect -46 130 -39 132
rect -33 132 -26 134
rect -33 130 -31 132
rect -29 130 -26 132
rect -46 125 -41 130
rect -33 128 -26 130
rect -31 125 -26 128
rect -24 125 -13 134
rect -11 125 -6 136
rect -4 134 3 136
rect -4 132 -1 134
rect 1 132 3 134
rect -4 130 3 132
rect 15 134 22 136
rect 15 132 17 134
rect 19 132 22 134
rect -4 125 1 130
rect 15 129 22 132
rect 24 141 33 143
rect 24 139 28 141
rect 30 139 33 141
rect 24 129 33 139
rect 26 123 33 129
rect 35 123 40 143
rect 42 136 47 143
rect 85 140 90 143
rect 75 137 80 140
rect 42 134 49 136
rect 42 132 45 134
rect 47 132 49 134
rect 42 130 49 132
rect 53 134 60 137
rect 53 132 55 134
rect 57 132 60 134
rect 42 123 47 130
rect 53 127 60 132
rect 53 125 55 127
rect 57 125 60 127
rect 53 123 60 125
rect 62 127 70 137
rect 62 125 65 127
rect 67 125 70 127
rect 62 123 70 125
rect 72 135 80 137
rect 72 133 75 135
rect 77 133 80 135
rect 72 130 80 133
rect 82 138 90 140
rect 82 136 85 138
rect 87 136 90 138
rect 82 130 90 136
rect 92 136 97 143
rect 141 144 147 146
rect 141 142 143 144
rect 145 142 147 144
rect 141 137 147 142
rect 92 134 99 136
rect 92 132 95 134
rect 97 132 99 134
rect 130 135 137 137
rect 130 133 132 135
rect 134 133 137 135
rect 92 130 99 132
rect 72 123 77 130
rect 108 129 113 132
rect 106 127 113 129
rect 106 125 108 127
rect 110 125 113 127
rect 106 123 113 125
rect 115 130 126 132
rect 130 131 137 133
rect 115 128 122 130
rect 124 128 126 130
rect 115 123 126 128
rect 132 125 137 131
rect 139 135 147 137
rect 195 144 201 146
rect 195 142 197 144
rect 199 142 201 144
rect 139 125 149 135
rect 141 123 149 125
rect 151 123 156 135
rect 158 127 166 135
rect 158 125 161 127
rect 163 125 166 127
rect 158 123 166 125
rect 168 133 176 135
rect 168 131 171 133
rect 173 131 176 133
rect 168 123 176 131
rect 178 133 186 135
rect 178 131 181 133
rect 183 131 186 133
rect 178 123 186 131
rect 195 129 203 142
rect 205 129 210 142
rect 212 134 220 142
rect 212 132 215 134
rect 217 132 220 134
rect 212 129 220 132
rect 222 137 227 142
rect 234 141 240 143
rect 234 139 236 141
rect 238 140 240 141
rect 257 144 263 146
rect 257 142 259 144
rect 261 142 263 144
rect 238 139 242 140
rect 234 137 242 139
rect 222 133 230 137
rect 222 131 225 133
rect 227 131 230 133
rect 222 129 230 131
rect 225 124 230 129
rect 232 129 242 137
rect 244 135 249 140
rect 244 133 251 135
rect 244 131 247 133
rect 249 131 251 133
rect 244 129 251 131
rect 257 129 265 142
rect 267 129 272 142
rect 274 134 282 142
rect 274 132 277 134
rect 279 132 282 134
rect 274 129 282 132
rect 284 137 289 142
rect 284 133 292 137
rect 284 131 287 133
rect 289 131 292 133
rect 284 129 292 131
rect 232 124 240 129
rect 287 124 292 129
rect 294 135 301 137
rect 294 133 297 135
rect 299 134 301 135
rect 359 144 365 146
rect 359 142 361 144
rect 363 142 365 144
rect 359 137 365 142
rect 299 133 303 134
rect 294 124 303 133
rect 298 123 303 124
rect 305 129 310 134
rect 348 135 355 137
rect 348 133 350 135
rect 352 133 355 135
rect 326 129 331 132
rect 305 127 312 129
rect 305 125 308 127
rect 310 125 312 127
rect 305 123 312 125
rect 324 127 331 129
rect 324 125 326 127
rect 328 125 331 127
rect 324 123 331 125
rect 333 130 344 132
rect 348 131 355 133
rect 333 128 340 130
rect 342 128 344 130
rect 333 123 344 128
rect 350 125 355 131
rect 357 135 365 137
rect 413 144 419 146
rect 413 142 415 144
rect 417 142 419 144
rect 357 125 367 135
rect 359 123 367 125
rect 369 123 374 135
rect 376 127 384 135
rect 376 125 379 127
rect 381 125 384 127
rect 376 123 384 125
rect 386 133 394 135
rect 386 131 389 133
rect 391 131 394 133
rect 386 123 394 131
rect 396 133 404 135
rect 396 131 399 133
rect 401 131 404 133
rect 396 123 404 131
rect 413 129 421 142
rect 423 129 428 142
rect 430 134 438 142
rect 430 132 433 134
rect 435 132 438 134
rect 430 129 438 132
rect 440 137 445 142
rect 452 141 458 143
rect 452 139 454 141
rect 456 140 458 141
rect 475 144 481 146
rect 475 142 477 144
rect 479 142 481 144
rect 456 139 460 140
rect 452 137 460 139
rect 440 133 448 137
rect 440 131 443 133
rect 445 131 448 133
rect 440 129 448 131
rect 443 124 448 129
rect 450 129 460 137
rect 462 135 467 140
rect 462 133 469 135
rect 462 131 465 133
rect 467 131 469 133
rect 462 129 469 131
rect 475 129 483 142
rect 485 129 490 142
rect 492 134 500 142
rect 492 132 495 134
rect 497 132 500 134
rect 492 129 500 132
rect 502 137 507 142
rect 502 133 510 137
rect 502 131 505 133
rect 507 131 510 133
rect 502 129 510 131
rect 450 124 458 129
rect 505 124 510 129
rect 512 135 519 137
rect 512 133 515 135
rect 517 134 519 135
rect 555 136 560 143
rect 553 134 560 136
rect 517 133 521 134
rect 512 124 521 133
rect 516 123 521 124
rect 523 129 528 134
rect 553 132 555 134
rect 557 132 560 134
rect 553 129 560 132
rect 562 141 571 143
rect 562 139 566 141
rect 568 139 571 141
rect 562 129 571 139
rect 523 127 530 129
rect 523 125 526 127
rect 528 125 530 127
rect 523 123 530 125
rect 564 123 571 129
rect 573 123 578 143
rect 580 136 585 143
rect 623 140 628 143
rect 613 137 618 140
rect 580 134 587 136
rect 580 132 583 134
rect 585 132 587 134
rect 580 130 587 132
rect 591 134 598 137
rect 591 132 593 134
rect 595 132 598 134
rect 580 123 585 130
rect 591 127 598 132
rect 591 125 593 127
rect 595 125 598 127
rect 591 123 598 125
rect 600 127 608 137
rect 600 125 603 127
rect 605 125 608 127
rect 600 123 608 125
rect 610 135 618 137
rect 610 133 613 135
rect 615 133 618 135
rect 610 130 618 133
rect 620 138 628 140
rect 620 136 623 138
rect 625 136 628 138
rect 620 130 628 136
rect 630 136 635 143
rect 630 134 637 136
rect 630 132 633 134
rect 635 132 637 134
rect 630 130 637 132
rect 610 123 615 130
rect -148 29 -141 31
rect -190 26 -185 29
rect -192 24 -185 26
rect -192 22 -190 24
rect -188 22 -185 24
rect -192 20 -185 22
rect -183 20 -172 29
rect -181 18 -172 20
rect -170 18 -165 29
rect -163 24 -158 29
rect -148 27 -146 29
rect -144 27 -141 29
rect -148 25 -141 27
rect -163 22 -156 24
rect -146 22 -141 25
rect -139 26 -128 31
rect -113 29 -105 31
rect -139 24 -132 26
rect -130 24 -128 26
rect -139 22 -128 24
rect -122 23 -117 29
rect -163 20 -160 22
rect -158 20 -156 22
rect -163 18 -156 20
rect -181 12 -174 18
rect -124 21 -117 23
rect -124 19 -122 21
rect -120 19 -117 21
rect -124 17 -117 19
rect -115 19 -105 29
rect -103 19 -98 31
rect -96 29 -88 31
rect -96 27 -93 29
rect -91 27 -88 29
rect -96 19 -88 27
rect -86 23 -78 31
rect -86 21 -83 23
rect -81 21 -78 23
rect -86 19 -78 21
rect -76 23 -68 31
rect -29 25 -24 30
rect -76 21 -73 23
rect -71 21 -68 23
rect -76 19 -68 21
rect -115 17 -107 19
rect -181 10 -179 12
rect -177 10 -174 12
rect -181 8 -174 10
rect -113 12 -107 17
rect -113 10 -111 12
rect -109 10 -107 12
rect -113 8 -107 10
rect -59 12 -51 25
rect -49 12 -44 25
rect -42 22 -34 25
rect -42 20 -39 22
rect -37 20 -34 22
rect -42 12 -34 20
rect -32 23 -24 25
rect -32 21 -29 23
rect -27 21 -24 23
rect -32 17 -24 21
rect -22 25 -14 30
rect 44 30 49 31
rect 33 25 38 30
rect -22 17 -12 25
rect -32 12 -27 17
rect -20 15 -12 17
rect -20 13 -18 15
rect -16 14 -12 15
rect -10 23 -3 25
rect -10 21 -7 23
rect -5 21 -3 23
rect -10 19 -3 21
rect -10 14 -5 19
rect -16 13 -14 14
rect -59 10 -57 12
rect -55 10 -53 12
rect -59 8 -53 10
rect -20 11 -14 13
rect 3 12 11 25
rect 13 12 18 25
rect 20 22 28 25
rect 20 20 23 22
rect 25 20 28 22
rect 20 12 28 20
rect 30 23 38 25
rect 30 21 33 23
rect 35 21 38 23
rect 30 17 38 21
rect 40 21 49 30
rect 40 19 43 21
rect 45 20 49 21
rect 51 29 58 31
rect 51 27 54 29
rect 56 27 58 29
rect 51 25 58 27
rect 70 29 77 31
rect 70 27 72 29
rect 74 27 77 29
rect 70 25 77 27
rect 51 20 56 25
rect 72 22 77 25
rect 79 26 90 31
rect 105 29 113 31
rect 79 24 86 26
rect 88 24 90 26
rect 79 22 90 24
rect 96 23 101 29
rect 45 19 47 20
rect 40 17 47 19
rect 30 12 35 17
rect 3 10 5 12
rect 7 10 9 12
rect 3 8 9 10
rect 94 21 101 23
rect 94 19 96 21
rect 98 19 101 21
rect 94 17 101 19
rect 103 19 113 29
rect 115 19 120 31
rect 122 29 130 31
rect 122 27 125 29
rect 127 27 130 29
rect 122 19 130 27
rect 132 23 140 31
rect 132 21 135 23
rect 137 21 140 23
rect 132 19 140 21
rect 142 23 150 31
rect 189 25 194 30
rect 142 21 145 23
rect 147 21 150 23
rect 142 19 150 21
rect 103 17 111 19
rect 105 12 111 17
rect 105 10 107 12
rect 109 10 111 12
rect 105 8 111 10
rect 159 12 167 25
rect 169 12 174 25
rect 176 22 184 25
rect 176 20 179 22
rect 181 20 184 22
rect 176 12 184 20
rect 186 23 194 25
rect 186 21 189 23
rect 191 21 194 23
rect 186 17 194 21
rect 196 25 204 30
rect 262 30 267 31
rect 251 25 256 30
rect 196 17 206 25
rect 186 12 191 17
rect 198 15 206 17
rect 198 13 200 15
rect 202 14 206 15
rect 208 23 215 25
rect 208 21 211 23
rect 213 21 215 23
rect 208 19 215 21
rect 208 14 213 19
rect 202 13 204 14
rect 159 10 161 12
rect 163 10 165 12
rect 159 8 165 10
rect 198 11 204 13
rect 221 12 229 25
rect 231 12 236 25
rect 238 22 246 25
rect 238 20 241 22
rect 243 20 246 22
rect 238 12 246 20
rect 248 23 256 25
rect 248 21 251 23
rect 253 21 256 23
rect 248 17 256 21
rect 258 21 267 30
rect 258 19 261 21
rect 263 20 267 21
rect 269 29 276 31
rect 269 27 272 29
rect 274 27 276 29
rect 269 25 276 27
rect 290 29 297 31
rect 290 27 292 29
rect 294 27 297 29
rect 290 25 297 27
rect 269 20 274 25
rect 292 22 297 25
rect 299 26 310 31
rect 325 29 333 31
rect 299 24 306 26
rect 308 24 310 26
rect 299 22 310 24
rect 316 23 321 29
rect 263 19 265 20
rect 258 17 265 19
rect 248 12 253 17
rect 221 10 223 12
rect 225 10 227 12
rect 221 8 227 10
rect 314 21 321 23
rect 314 19 316 21
rect 318 19 321 21
rect 314 17 321 19
rect 323 19 333 29
rect 335 19 340 31
rect 342 29 350 31
rect 342 27 345 29
rect 347 27 350 29
rect 342 19 350 27
rect 352 23 360 31
rect 352 21 355 23
rect 357 21 360 23
rect 352 19 360 21
rect 362 23 370 31
rect 409 25 414 30
rect 362 21 365 23
rect 367 21 370 23
rect 362 19 370 21
rect 323 17 331 19
rect 325 12 331 17
rect 325 10 327 12
rect 329 10 331 12
rect 325 8 331 10
rect 379 12 387 25
rect 389 12 394 25
rect 396 22 404 25
rect 396 20 399 22
rect 401 20 404 22
rect 396 12 404 20
rect 406 23 414 25
rect 406 21 409 23
rect 411 21 414 23
rect 406 17 414 21
rect 416 25 424 30
rect 482 30 487 31
rect 471 25 476 30
rect 416 17 426 25
rect 406 12 411 17
rect 418 15 426 17
rect 418 13 420 15
rect 422 14 426 15
rect 428 23 435 25
rect 428 21 431 23
rect 433 21 435 23
rect 428 19 435 21
rect 428 14 433 19
rect 422 13 424 14
rect 379 10 381 12
rect 383 10 385 12
rect 379 8 385 10
rect 418 11 424 13
rect 441 12 449 25
rect 451 12 456 25
rect 458 22 466 25
rect 458 20 461 22
rect 463 20 466 22
rect 458 12 466 20
rect 468 23 476 25
rect 468 21 471 23
rect 473 21 476 23
rect 468 17 476 21
rect 478 21 487 30
rect 478 19 481 21
rect 483 20 487 21
rect 489 29 496 31
rect 489 27 492 29
rect 494 27 496 29
rect 489 25 496 27
rect 523 25 530 31
rect 489 20 494 25
rect 512 22 519 25
rect 512 20 514 22
rect 516 20 519 22
rect 483 19 485 20
rect 478 17 485 19
rect 468 12 473 17
rect 441 10 443 12
rect 445 10 447 12
rect 441 8 447 10
rect 512 18 519 20
rect 514 11 519 18
rect 521 15 530 25
rect 521 13 525 15
rect 527 13 530 15
rect 521 11 530 13
rect 532 11 537 31
rect 539 24 544 31
rect 550 29 557 31
rect 550 27 552 29
rect 554 27 557 29
rect 539 22 546 24
rect 539 20 542 22
rect 544 20 546 22
rect 539 18 546 20
rect 550 22 557 27
rect 550 20 552 22
rect 554 20 557 22
rect 539 11 544 18
rect 550 17 557 20
rect 559 29 567 31
rect 559 27 562 29
rect 564 27 567 29
rect 559 17 567 27
rect 569 24 574 31
rect 569 21 577 24
rect 569 19 572 21
rect 574 19 577 21
rect 569 17 577 19
rect 572 14 577 17
rect 579 18 587 24
rect 579 16 582 18
rect 584 16 587 18
rect 579 14 587 16
rect 582 11 587 14
rect 589 22 596 24
rect 589 20 592 22
rect 594 20 596 22
rect 589 18 596 20
rect 589 11 594 18
rect -175 0 -169 2
rect -175 -2 -173 0
rect -171 -2 -169 0
rect -175 -7 -169 -2
rect -186 -9 -179 -7
rect -186 -11 -184 -9
rect -182 -11 -179 -9
rect -208 -15 -203 -12
rect -210 -17 -203 -15
rect -210 -19 -208 -17
rect -206 -19 -203 -17
rect -210 -21 -203 -19
rect -201 -14 -190 -12
rect -186 -13 -179 -11
rect -201 -16 -194 -14
rect -192 -16 -190 -14
rect -201 -21 -190 -16
rect -184 -19 -179 -13
rect -177 -9 -169 -7
rect -121 0 -115 2
rect -121 -2 -119 0
rect -117 -2 -115 0
rect -177 -19 -167 -9
rect -175 -21 -167 -19
rect -165 -21 -160 -9
rect -158 -17 -150 -9
rect -158 -19 -155 -17
rect -153 -19 -150 -17
rect -158 -21 -150 -19
rect -148 -11 -140 -9
rect -148 -13 -145 -11
rect -143 -13 -140 -11
rect -148 -21 -140 -13
rect -138 -11 -130 -9
rect -138 -13 -135 -11
rect -133 -13 -130 -11
rect -138 -21 -130 -13
rect -121 -15 -113 -2
rect -111 -15 -106 -2
rect -104 -10 -96 -2
rect -104 -12 -101 -10
rect -99 -12 -96 -10
rect -104 -15 -96 -12
rect -94 -7 -89 -2
rect -82 -3 -76 -1
rect -82 -5 -80 -3
rect -78 -4 -76 -3
rect -59 0 -53 2
rect -59 -2 -57 0
rect -55 -2 -53 0
rect -78 -5 -74 -4
rect -82 -7 -74 -5
rect -94 -11 -86 -7
rect -94 -13 -91 -11
rect -89 -13 -86 -11
rect -94 -15 -86 -13
rect -91 -20 -86 -15
rect -84 -15 -74 -7
rect -72 -9 -67 -4
rect -72 -11 -65 -9
rect -72 -13 -69 -11
rect -67 -13 -65 -11
rect -72 -15 -65 -13
rect -59 -15 -51 -2
rect -49 -15 -44 -2
rect -42 -10 -34 -2
rect -42 -12 -39 -10
rect -37 -12 -34 -10
rect -42 -15 -34 -12
rect -32 -7 -27 -2
rect -32 -11 -24 -7
rect -32 -13 -29 -11
rect -27 -13 -24 -11
rect -32 -15 -24 -13
rect -84 -20 -76 -15
rect -29 -20 -24 -15
rect -22 -9 -15 -7
rect -22 -11 -19 -9
rect -17 -10 -15 -9
rect 45 0 51 2
rect 45 -2 47 0
rect 49 -2 51 0
rect 45 -7 51 -2
rect -17 -11 -13 -10
rect -22 -20 -13 -11
rect -18 -21 -13 -20
rect -11 -15 -6 -10
rect 34 -9 41 -7
rect 34 -11 36 -9
rect 38 -11 41 -9
rect 12 -15 17 -12
rect -11 -17 -4 -15
rect -11 -19 -8 -17
rect -6 -19 -4 -17
rect -11 -21 -4 -19
rect 10 -17 17 -15
rect 10 -19 12 -17
rect 14 -19 17 -17
rect 10 -21 17 -19
rect 19 -14 30 -12
rect 34 -13 41 -11
rect 19 -16 26 -14
rect 28 -16 30 -14
rect 19 -21 30 -16
rect 36 -19 41 -13
rect 43 -9 51 -7
rect 99 0 105 2
rect 99 -2 101 0
rect 103 -2 105 0
rect 43 -19 53 -9
rect 45 -21 53 -19
rect 55 -21 60 -9
rect 62 -17 70 -9
rect 62 -19 65 -17
rect 67 -19 70 -17
rect 62 -21 70 -19
rect 72 -11 80 -9
rect 72 -13 75 -11
rect 77 -13 80 -11
rect 72 -21 80 -13
rect 82 -11 90 -9
rect 82 -13 85 -11
rect 87 -13 90 -11
rect 82 -21 90 -13
rect 99 -15 107 -2
rect 109 -15 114 -2
rect 116 -10 124 -2
rect 116 -12 119 -10
rect 121 -12 124 -10
rect 116 -15 124 -12
rect 126 -7 131 -2
rect 138 -3 144 -1
rect 138 -5 140 -3
rect 142 -4 144 -3
rect 161 0 167 2
rect 161 -2 163 0
rect 165 -2 167 0
rect 142 -5 146 -4
rect 138 -7 146 -5
rect 126 -11 134 -7
rect 126 -13 129 -11
rect 131 -13 134 -11
rect 126 -15 134 -13
rect 129 -20 134 -15
rect 136 -15 146 -7
rect 148 -9 153 -4
rect 148 -11 155 -9
rect 148 -13 151 -11
rect 153 -13 155 -11
rect 148 -15 155 -13
rect 161 -15 169 -2
rect 171 -15 176 -2
rect 178 -10 186 -2
rect 178 -12 181 -10
rect 183 -12 186 -10
rect 178 -15 186 -12
rect 188 -7 193 -2
rect 188 -11 196 -7
rect 188 -13 191 -11
rect 193 -13 196 -11
rect 188 -15 196 -13
rect 136 -20 144 -15
rect 191 -20 196 -15
rect 198 -9 205 -7
rect 198 -11 201 -9
rect 203 -10 205 -9
rect 262 0 268 2
rect 262 -2 264 0
rect 266 -2 268 0
rect 262 -7 268 -2
rect 203 -11 207 -10
rect 198 -20 207 -11
rect 202 -21 207 -20
rect 209 -15 214 -10
rect 251 -9 258 -7
rect 251 -11 253 -9
rect 255 -11 258 -9
rect 229 -15 234 -12
rect 209 -17 216 -15
rect 209 -19 212 -17
rect 214 -19 216 -17
rect 209 -21 216 -19
rect 227 -17 234 -15
rect 227 -19 229 -17
rect 231 -19 234 -17
rect 227 -21 234 -19
rect 236 -14 247 -12
rect 251 -13 258 -11
rect 236 -16 243 -14
rect 245 -16 247 -14
rect 236 -21 247 -16
rect 253 -19 258 -13
rect 260 -9 268 -7
rect 316 0 322 2
rect 316 -2 318 0
rect 320 -2 322 0
rect 260 -19 270 -9
rect 262 -21 270 -19
rect 272 -21 277 -9
rect 279 -17 287 -9
rect 279 -19 282 -17
rect 284 -19 287 -17
rect 279 -21 287 -19
rect 289 -11 297 -9
rect 289 -13 292 -11
rect 294 -13 297 -11
rect 289 -21 297 -13
rect 299 -11 307 -9
rect 299 -13 302 -11
rect 304 -13 307 -11
rect 299 -21 307 -13
rect 316 -15 324 -2
rect 326 -15 331 -2
rect 333 -10 341 -2
rect 333 -12 336 -10
rect 338 -12 341 -10
rect 333 -15 341 -12
rect 343 -7 348 -2
rect 355 -3 361 -1
rect 355 -5 357 -3
rect 359 -4 361 -3
rect 378 0 384 2
rect 378 -2 380 0
rect 382 -2 384 0
rect 359 -5 363 -4
rect 355 -7 363 -5
rect 343 -11 351 -7
rect 343 -13 346 -11
rect 348 -13 351 -11
rect 343 -15 351 -13
rect 346 -20 351 -15
rect 353 -15 363 -7
rect 365 -9 370 -4
rect 365 -11 372 -9
rect 365 -13 368 -11
rect 370 -13 372 -11
rect 365 -15 372 -13
rect 378 -15 386 -2
rect 388 -15 393 -2
rect 395 -10 403 -2
rect 395 -12 398 -10
rect 400 -12 403 -10
rect 395 -15 403 -12
rect 405 -7 410 -2
rect 405 -11 413 -7
rect 405 -13 408 -11
rect 410 -13 413 -11
rect 405 -15 413 -13
rect 353 -20 361 -15
rect 408 -20 413 -15
rect 415 -9 422 -7
rect 415 -11 418 -9
rect 420 -10 422 -9
rect 457 -8 462 -1
rect 455 -10 462 -8
rect 420 -11 424 -10
rect 415 -20 424 -11
rect 419 -21 424 -20
rect 426 -15 431 -10
rect 455 -12 457 -10
rect 459 -12 462 -10
rect 455 -15 462 -12
rect 464 -3 473 -1
rect 464 -5 468 -3
rect 470 -5 473 -3
rect 464 -15 473 -5
rect 426 -17 433 -15
rect 426 -19 429 -17
rect 431 -19 433 -17
rect 426 -21 433 -19
rect 466 -21 473 -15
rect 475 -21 480 -1
rect 482 -8 487 -1
rect 525 -4 530 -1
rect 515 -7 520 -4
rect 482 -10 489 -8
rect 482 -12 485 -10
rect 487 -12 489 -10
rect 482 -14 489 -12
rect 493 -10 500 -7
rect 493 -12 495 -10
rect 497 -12 500 -10
rect 482 -21 487 -14
rect 493 -17 500 -12
rect 493 -19 495 -17
rect 497 -19 500 -17
rect 493 -21 500 -19
rect 502 -17 510 -7
rect 502 -19 505 -17
rect 507 -19 510 -17
rect 502 -21 510 -19
rect 512 -9 520 -7
rect 512 -11 515 -9
rect 517 -11 520 -9
rect 512 -14 520 -11
rect 522 -6 530 -4
rect 522 -8 525 -6
rect 527 -8 530 -6
rect 522 -14 530 -8
rect 532 -8 537 -1
rect 532 -10 539 -8
rect 532 -12 535 -10
rect 537 -12 539 -10
rect 532 -14 539 -12
rect 512 -21 517 -14
<< pdif >>
rect 53 205 59 207
rect 44 200 49 205
rect 42 198 49 200
rect 42 196 44 198
rect 46 196 49 198
rect 42 191 49 196
rect 42 189 44 191
rect 46 189 49 191
rect 42 187 49 189
rect 51 203 59 205
rect 51 201 54 203
rect 56 201 59 203
rect 51 194 59 201
rect 61 205 69 207
rect 61 203 64 205
rect 66 203 69 205
rect 61 198 69 203
rect 61 196 64 198
rect 66 196 69 198
rect 61 194 69 196
rect 71 205 78 207
rect 93 205 99 207
rect 71 203 74 205
rect 76 203 78 205
rect 71 194 78 203
rect 84 200 89 205
rect 82 198 89 200
rect 82 196 84 198
rect 86 196 89 198
rect 51 187 57 194
rect 82 191 89 196
rect 82 189 84 191
rect 86 189 89 191
rect 82 187 89 189
rect 91 203 99 205
rect 91 201 94 203
rect 96 201 99 203
rect 91 194 99 201
rect 101 205 109 207
rect 101 203 104 205
rect 106 203 109 205
rect 101 198 109 203
rect 101 196 104 198
rect 106 196 109 198
rect 101 194 109 196
rect 111 205 118 207
rect 136 205 142 207
rect 111 203 114 205
rect 116 203 118 205
rect 111 194 118 203
rect 127 200 132 205
rect 125 198 132 200
rect 125 196 127 198
rect 129 196 132 198
rect 91 187 97 194
rect 125 191 132 196
rect 125 189 127 191
rect 129 189 132 191
rect 125 187 132 189
rect 134 203 142 205
rect 134 201 137 203
rect 139 201 142 203
rect 134 194 142 201
rect 144 205 152 207
rect 144 203 147 205
rect 149 203 152 205
rect 144 198 152 203
rect 144 196 147 198
rect 149 196 152 198
rect 144 194 152 196
rect 154 205 161 207
rect 240 205 246 207
rect 154 203 157 205
rect 159 203 161 205
rect 154 194 161 203
rect 231 200 236 205
rect 229 198 236 200
rect 229 196 231 198
rect 233 196 236 198
rect 134 187 140 194
rect 229 191 236 196
rect 229 189 231 191
rect 233 189 236 191
rect 229 187 236 189
rect 238 203 246 205
rect 238 201 241 203
rect 243 201 246 203
rect 238 194 246 201
rect 248 205 256 207
rect 248 203 251 205
rect 253 203 256 205
rect 248 198 256 203
rect 248 196 251 198
rect 253 196 256 198
rect 248 194 256 196
rect 258 205 265 207
rect 282 205 288 207
rect 258 203 261 205
rect 263 203 265 205
rect 258 194 265 203
rect 273 200 278 205
rect 271 198 278 200
rect 271 196 273 198
rect 275 196 278 198
rect 238 187 244 194
rect 271 191 278 196
rect 271 189 273 191
rect 275 189 278 191
rect 271 187 278 189
rect 280 203 288 205
rect 280 201 283 203
rect 285 201 288 203
rect 280 194 288 201
rect 290 205 298 207
rect 290 203 293 205
rect 295 203 298 205
rect 290 198 298 203
rect 290 196 293 198
rect 295 196 298 198
rect 290 194 298 196
rect 300 205 307 207
rect 326 205 332 207
rect 300 203 303 205
rect 305 203 307 205
rect 300 194 307 203
rect 317 200 322 205
rect 315 198 322 200
rect 315 196 317 198
rect 319 196 322 198
rect 280 187 286 194
rect 315 191 322 196
rect 315 189 317 191
rect 319 189 322 191
rect 315 187 322 189
rect 324 203 332 205
rect 324 201 327 203
rect 329 201 332 203
rect 324 194 332 201
rect 334 205 342 207
rect 334 203 337 205
rect 339 203 342 205
rect 334 198 342 203
rect 334 196 337 198
rect 339 196 342 198
rect 334 194 342 196
rect 344 205 351 207
rect 395 205 401 207
rect 344 203 347 205
rect 349 203 351 205
rect 344 194 351 203
rect 386 200 391 205
rect 384 198 391 200
rect 384 196 386 198
rect 388 196 391 198
rect 324 187 330 194
rect 384 191 391 196
rect 384 189 386 191
rect 388 189 391 191
rect 384 187 391 189
rect 393 203 401 205
rect 393 201 396 203
rect 398 201 401 203
rect 393 194 401 201
rect 403 205 411 207
rect 403 203 406 205
rect 408 203 411 205
rect 403 198 411 203
rect 403 196 406 198
rect 408 196 411 198
rect 403 194 411 196
rect 413 205 420 207
rect 439 205 445 207
rect 413 203 416 205
rect 418 203 420 205
rect 413 194 420 203
rect 430 200 435 205
rect 428 198 435 200
rect 428 196 430 198
rect 432 196 435 198
rect 393 187 399 194
rect 428 191 435 196
rect 428 189 430 191
rect 432 189 435 191
rect 428 187 435 189
rect 437 203 445 205
rect 437 201 440 203
rect 442 201 445 203
rect 437 194 445 201
rect 447 205 455 207
rect 447 203 450 205
rect 452 203 455 205
rect 447 198 455 203
rect 447 196 450 198
rect 452 196 455 198
rect 447 194 455 196
rect 457 205 464 207
rect 481 205 487 207
rect 457 203 460 205
rect 462 203 464 205
rect 457 194 464 203
rect 472 200 477 205
rect 470 198 477 200
rect 470 196 472 198
rect 474 196 477 198
rect 437 187 443 194
rect 470 191 477 196
rect 470 189 472 191
rect 474 189 477 191
rect 470 187 477 189
rect 479 203 487 205
rect 479 201 482 203
rect 484 201 487 203
rect 479 194 487 201
rect 489 205 497 207
rect 489 203 492 205
rect 494 203 497 205
rect 489 198 497 203
rect 489 196 492 198
rect 494 196 497 198
rect 489 194 497 196
rect 499 205 506 207
rect 522 205 528 207
rect 499 203 502 205
rect 504 203 506 205
rect 499 194 506 203
rect 513 200 518 205
rect 511 198 518 200
rect 511 196 513 198
rect 515 196 518 198
rect 479 187 485 194
rect 511 191 518 196
rect 511 189 513 191
rect 515 189 518 191
rect 511 187 518 189
rect 520 203 528 205
rect 520 201 523 203
rect 525 201 528 203
rect 520 194 528 201
rect 530 205 538 207
rect 530 203 533 205
rect 535 203 538 205
rect 530 198 538 203
rect 530 196 533 198
rect 535 196 538 198
rect 530 194 538 196
rect 540 205 547 207
rect 565 205 571 207
rect 540 203 543 205
rect 545 203 547 205
rect 540 194 547 203
rect 556 200 561 205
rect 554 198 561 200
rect 554 196 556 198
rect 558 196 561 198
rect 520 187 526 194
rect 554 191 561 196
rect 554 189 556 191
rect 558 189 561 191
rect 554 187 561 189
rect 563 203 571 205
rect 563 201 566 203
rect 568 201 571 203
rect 563 194 571 201
rect 573 205 581 207
rect 573 203 576 205
rect 578 203 581 205
rect 573 198 581 203
rect 573 196 576 198
rect 578 196 581 198
rect 573 194 581 196
rect 583 205 590 207
rect 605 205 611 207
rect 583 203 586 205
rect 588 203 590 205
rect 583 194 590 203
rect 596 200 601 205
rect 594 198 601 200
rect 594 196 596 198
rect 598 196 601 198
rect 563 187 569 194
rect 594 191 601 196
rect 594 189 596 191
rect 598 189 601 191
rect 594 187 601 189
rect 603 203 611 205
rect 603 201 606 203
rect 608 201 611 203
rect 603 194 611 201
rect 613 205 621 207
rect 613 203 616 205
rect 618 203 621 205
rect 613 198 621 203
rect 613 196 616 198
rect 618 196 621 198
rect 613 194 621 196
rect 623 205 630 207
rect 648 205 654 207
rect 623 203 626 205
rect 628 203 630 205
rect 623 194 630 203
rect 639 200 644 205
rect 637 198 644 200
rect 637 196 639 198
rect 641 196 644 198
rect 603 187 609 194
rect 637 191 644 196
rect 637 189 639 191
rect 641 189 644 191
rect 637 187 644 189
rect 646 203 654 205
rect 646 201 649 203
rect 651 201 654 203
rect 646 194 654 201
rect 656 205 664 207
rect 656 203 659 205
rect 661 203 664 205
rect 656 198 664 203
rect 656 196 659 198
rect 661 196 664 198
rect 656 194 664 196
rect 666 205 673 207
rect 666 203 669 205
rect 671 203 673 205
rect 666 194 673 203
rect 646 187 652 194
rect -75 108 -68 110
rect -75 106 -73 108
rect -71 106 -68 108
rect -75 101 -68 106
rect -75 99 -73 101
rect -71 99 -68 101
rect -75 97 -68 99
rect -73 92 -68 97
rect -66 103 -60 110
rect -33 108 -26 110
rect -33 106 -31 108
rect -29 106 -26 108
rect -66 96 -58 103
rect -66 94 -63 96
rect -61 94 -58 96
rect -66 92 -58 94
rect -64 90 -58 92
rect -56 101 -48 103
rect -56 99 -53 101
rect -51 99 -48 101
rect -56 94 -48 99
rect -56 92 -53 94
rect -51 92 -48 94
rect -56 90 -48 92
rect -46 94 -39 103
rect -33 101 -26 106
rect -33 99 -31 101
rect -29 99 -26 101
rect -33 97 -26 99
rect -46 92 -43 94
rect -41 92 -39 94
rect -31 92 -26 97
rect -24 103 -18 110
rect 15 109 22 111
rect 15 107 17 109
rect 19 107 22 109
rect -24 96 -16 103
rect -24 94 -21 96
rect -19 94 -16 96
rect -24 92 -16 94
rect -46 90 -39 92
rect -22 90 -16 92
rect -14 101 -6 103
rect -14 99 -11 101
rect -9 99 -6 101
rect -14 94 -6 99
rect -14 92 -11 94
rect -9 92 -6 94
rect -14 90 -6 92
rect -4 94 3 103
rect 15 102 22 107
rect 15 100 17 102
rect 19 100 22 102
rect 15 98 22 100
rect -4 92 -1 94
rect 1 92 3 94
rect -4 90 3 92
rect 17 83 22 98
rect 24 94 32 111
rect 24 92 27 94
rect 29 92 32 94
rect 24 87 32 92
rect 24 85 27 87
rect 29 85 32 87
rect 24 83 32 85
rect 34 102 42 111
rect 34 100 37 102
rect 39 100 42 102
rect 34 95 42 100
rect 34 93 37 95
rect 39 93 42 95
rect 34 83 42 93
rect 44 94 60 111
rect 44 92 49 94
rect 51 92 60 94
rect 44 87 60 92
rect 44 85 49 87
rect 51 86 60 87
rect 62 86 67 111
rect 69 108 74 111
rect 106 109 113 111
rect 69 106 77 108
rect 69 104 72 106
rect 74 104 77 106
rect 69 95 77 104
rect 79 95 90 108
rect 69 86 74 95
rect 81 87 90 95
rect 51 85 58 86
rect 44 83 58 85
rect 81 85 84 87
rect 86 85 90 87
rect 81 83 90 85
rect 92 106 99 108
rect 92 104 95 106
rect 97 104 99 106
rect 92 99 99 104
rect 92 97 95 99
rect 97 97 99 99
rect 106 107 108 109
rect 110 107 113 109
rect 106 102 113 107
rect 106 100 108 102
rect 110 100 113 102
rect 106 98 113 100
rect 92 95 99 97
rect 92 83 97 95
rect 108 93 113 98
rect 115 94 124 111
rect 135 103 140 111
rect 115 93 119 94
rect 117 92 119 93
rect 121 92 124 94
rect 117 90 124 92
rect 133 101 140 103
rect 133 99 135 101
rect 137 99 140 101
rect 133 94 140 99
rect 133 92 135 94
rect 137 92 140 94
rect 133 90 140 92
rect 135 84 140 90
rect 142 95 150 111
rect 142 93 145 95
rect 147 93 150 95
rect 142 88 150 93
rect 142 86 145 88
rect 147 86 150 88
rect 142 84 150 86
rect 152 84 157 111
rect 159 109 167 111
rect 159 107 162 109
rect 164 107 167 109
rect 159 102 167 107
rect 159 100 162 102
rect 164 100 167 102
rect 159 84 167 100
rect 169 93 177 111
rect 169 91 172 93
rect 174 91 177 93
rect 169 84 177 91
rect 179 96 186 111
rect 197 96 202 111
rect 179 94 182 96
rect 184 94 186 96
rect 179 88 186 94
rect 195 94 202 96
rect 195 92 197 94
rect 199 92 202 94
rect 195 90 202 92
rect 179 86 182 88
rect 184 86 186 88
rect 179 84 186 86
rect 197 83 202 90
rect 204 102 212 111
rect 204 100 207 102
rect 209 100 212 102
rect 204 83 212 100
rect 214 109 222 111
rect 214 107 217 109
rect 219 107 222 109
rect 214 102 222 107
rect 214 100 217 102
rect 219 100 222 102
rect 214 83 222 100
rect 224 97 230 111
rect 224 87 232 97
rect 224 85 227 87
rect 229 85 232 87
rect 224 83 232 85
rect 234 94 242 97
rect 234 92 237 94
rect 239 92 242 94
rect 234 83 242 92
rect 244 94 251 97
rect 257 96 262 111
rect 244 92 247 94
rect 249 92 251 94
rect 244 87 251 92
rect 255 94 262 96
rect 255 92 257 94
rect 259 92 262 94
rect 255 90 262 92
rect 244 85 247 87
rect 249 85 251 87
rect 244 83 251 85
rect 257 83 262 90
rect 264 102 272 111
rect 264 100 267 102
rect 269 100 272 102
rect 264 83 272 100
rect 274 109 282 111
rect 274 107 277 109
rect 279 107 282 109
rect 274 102 282 107
rect 274 100 277 102
rect 279 100 282 102
rect 274 83 282 100
rect 284 104 291 111
rect 324 109 331 111
rect 324 107 326 109
rect 328 107 331 109
rect 284 90 293 104
rect 295 102 303 104
rect 295 100 298 102
rect 300 100 303 102
rect 295 90 303 100
rect 305 94 313 104
rect 324 102 331 107
rect 324 100 326 102
rect 328 100 331 102
rect 324 98 331 100
rect 305 92 308 94
rect 310 92 313 94
rect 326 93 331 98
rect 333 94 342 111
rect 353 103 358 111
rect 333 93 337 94
rect 305 90 313 92
rect 284 87 291 90
rect 284 85 287 87
rect 289 85 291 87
rect 335 92 337 93
rect 339 92 342 94
rect 335 90 342 92
rect 351 101 358 103
rect 351 99 353 101
rect 355 99 358 101
rect 351 94 358 99
rect 351 92 353 94
rect 355 92 358 94
rect 351 90 358 92
rect 284 83 291 85
rect 353 84 358 90
rect 360 95 368 111
rect 360 93 363 95
rect 365 93 368 95
rect 360 88 368 93
rect 360 86 363 88
rect 365 86 368 88
rect 360 84 368 86
rect 370 84 375 111
rect 377 109 385 111
rect 377 107 380 109
rect 382 107 385 109
rect 377 102 385 107
rect 377 100 380 102
rect 382 100 385 102
rect 377 84 385 100
rect 387 93 395 111
rect 387 91 390 93
rect 392 91 395 93
rect 387 84 395 91
rect 397 96 404 111
rect 415 96 420 111
rect 397 94 400 96
rect 402 94 404 96
rect 397 88 404 94
rect 413 94 420 96
rect 413 92 415 94
rect 417 92 420 94
rect 413 90 420 92
rect 397 86 400 88
rect 402 86 404 88
rect 397 84 404 86
rect 415 83 420 90
rect 422 102 430 111
rect 422 100 425 102
rect 427 100 430 102
rect 422 83 430 100
rect 432 109 440 111
rect 432 107 435 109
rect 437 107 440 109
rect 432 102 440 107
rect 432 100 435 102
rect 437 100 440 102
rect 432 83 440 100
rect 442 97 448 111
rect 442 87 450 97
rect 442 85 445 87
rect 447 85 450 87
rect 442 83 450 85
rect 452 94 460 97
rect 452 92 455 94
rect 457 92 460 94
rect 452 83 460 92
rect 462 94 469 97
rect 475 96 480 111
rect 462 92 465 94
rect 467 92 469 94
rect 462 87 469 92
rect 473 94 480 96
rect 473 92 475 94
rect 477 92 480 94
rect 473 90 480 92
rect 462 85 465 87
rect 467 85 469 87
rect 462 83 469 85
rect 475 83 480 90
rect 482 102 490 111
rect 482 100 485 102
rect 487 100 490 102
rect 482 83 490 100
rect 492 109 500 111
rect 492 107 495 109
rect 497 107 500 109
rect 492 102 500 107
rect 492 100 495 102
rect 497 100 500 102
rect 492 83 500 100
rect 502 104 509 111
rect 553 109 560 111
rect 553 107 555 109
rect 557 107 560 109
rect 502 90 511 104
rect 513 102 521 104
rect 513 100 516 102
rect 518 100 521 102
rect 513 90 521 100
rect 523 94 531 104
rect 553 102 560 107
rect 553 100 555 102
rect 557 100 560 102
rect 553 98 560 100
rect 523 92 526 94
rect 528 92 531 94
rect 523 90 531 92
rect 502 87 509 90
rect 502 85 505 87
rect 507 85 509 87
rect 502 83 509 85
rect 555 83 560 98
rect 562 94 570 111
rect 562 92 565 94
rect 567 92 570 94
rect 562 87 570 92
rect 562 85 565 87
rect 567 85 570 87
rect 562 83 570 85
rect 572 102 580 111
rect 572 100 575 102
rect 577 100 580 102
rect 572 95 580 100
rect 572 93 575 95
rect 577 93 580 95
rect 572 83 580 93
rect 582 94 598 111
rect 582 92 587 94
rect 589 92 598 94
rect 582 87 598 92
rect 582 85 587 87
rect 589 86 598 87
rect 600 86 605 111
rect 607 108 612 111
rect 607 106 615 108
rect 607 104 610 106
rect 612 104 615 106
rect 607 95 615 104
rect 617 95 628 108
rect 607 86 612 95
rect 619 87 628 95
rect 589 85 596 86
rect 582 83 596 85
rect 619 85 622 87
rect 624 85 628 87
rect 619 83 628 85
rect 630 106 637 108
rect 630 104 633 106
rect 635 104 637 106
rect 630 99 637 104
rect 630 97 633 99
rect 635 97 637 99
rect 630 95 637 97
rect 630 83 635 95
rect -181 62 -175 64
rect -190 57 -185 62
rect -192 55 -185 57
rect -192 53 -190 55
rect -188 53 -185 55
rect -192 48 -185 53
rect -192 46 -190 48
rect -188 46 -185 48
rect -192 44 -185 46
rect -183 60 -175 62
rect -183 58 -180 60
rect -178 58 -175 60
rect -183 51 -175 58
rect -173 62 -165 64
rect -173 60 -170 62
rect -168 60 -165 62
rect -173 55 -165 60
rect -173 53 -170 55
rect -168 53 -165 55
rect -173 51 -165 53
rect -163 62 -156 64
rect -163 60 -160 62
rect -158 60 -156 62
rect -119 64 -114 70
rect -137 62 -130 64
rect -137 61 -135 62
rect -163 51 -156 60
rect -146 56 -141 61
rect -148 54 -141 56
rect -148 52 -146 54
rect -144 52 -141 54
rect -183 44 -177 51
rect -148 47 -141 52
rect -148 45 -146 47
rect -144 45 -141 47
rect -148 43 -141 45
rect -139 60 -135 61
rect -133 60 -130 62
rect -139 43 -130 60
rect -121 62 -114 64
rect -121 60 -119 62
rect -117 60 -114 62
rect -121 55 -114 60
rect -121 53 -119 55
rect -117 53 -114 55
rect -121 51 -114 53
rect -119 43 -114 51
rect -112 68 -104 70
rect -112 66 -109 68
rect -107 66 -104 68
rect -112 61 -104 66
rect -112 59 -109 61
rect -107 59 -104 61
rect -112 43 -104 59
rect -102 43 -97 70
rect -95 54 -87 70
rect -95 52 -92 54
rect -90 52 -87 54
rect -95 47 -87 52
rect -95 45 -92 47
rect -90 45 -87 47
rect -95 43 -87 45
rect -85 63 -77 70
rect -85 61 -82 63
rect -80 61 -77 63
rect -85 43 -77 61
rect -75 68 -68 70
rect -75 66 -72 68
rect -70 66 -68 68
rect -75 60 -68 66
rect -57 64 -52 71
rect -75 58 -72 60
rect -70 58 -68 60
rect -59 62 -52 64
rect -59 60 -57 62
rect -55 60 -52 62
rect -59 58 -52 60
rect -75 43 -68 58
rect -57 43 -52 58
rect -50 54 -42 71
rect -50 52 -47 54
rect -45 52 -42 54
rect -50 43 -42 52
rect -40 54 -32 71
rect -40 52 -37 54
rect -35 52 -32 54
rect -40 47 -32 52
rect -40 45 -37 47
rect -35 45 -32 47
rect -40 43 -32 45
rect -30 69 -22 71
rect -30 67 -27 69
rect -25 67 -22 69
rect -30 57 -22 67
rect -20 62 -12 71
rect -20 60 -17 62
rect -15 60 -12 62
rect -20 57 -12 60
rect -10 69 -3 71
rect -10 67 -7 69
rect -5 67 -3 69
rect -10 62 -3 67
rect 3 64 8 71
rect -10 60 -7 62
rect -5 60 -3 62
rect -10 57 -3 60
rect 1 62 8 64
rect 1 60 3 62
rect 5 60 8 62
rect 1 58 8 60
rect -30 43 -24 57
rect 3 43 8 58
rect 10 54 18 71
rect 10 52 13 54
rect 15 52 18 54
rect 10 43 18 52
rect 20 54 28 71
rect 20 52 23 54
rect 25 52 28 54
rect 20 47 28 52
rect 20 45 23 47
rect 25 45 28 47
rect 20 43 28 45
rect 30 69 37 71
rect 30 67 33 69
rect 35 67 37 69
rect 30 64 37 67
rect 30 50 39 64
rect 41 54 49 64
rect 41 52 44 54
rect 46 52 49 54
rect 41 50 49 52
rect 51 62 59 64
rect 51 60 54 62
rect 56 60 59 62
rect 99 64 104 70
rect 81 62 88 64
rect 81 61 83 62
rect 51 50 59 60
rect 72 56 77 61
rect 70 54 77 56
rect 70 52 72 54
rect 74 52 77 54
rect 30 43 37 50
rect 70 47 77 52
rect 70 45 72 47
rect 74 45 77 47
rect 70 43 77 45
rect 79 60 83 61
rect 85 60 88 62
rect 79 43 88 60
rect 97 62 104 64
rect 97 60 99 62
rect 101 60 104 62
rect 97 55 104 60
rect 97 53 99 55
rect 101 53 104 55
rect 97 51 104 53
rect 99 43 104 51
rect 106 68 114 70
rect 106 66 109 68
rect 111 66 114 68
rect 106 61 114 66
rect 106 59 109 61
rect 111 59 114 61
rect 106 43 114 59
rect 116 43 121 70
rect 123 54 131 70
rect 123 52 126 54
rect 128 52 131 54
rect 123 47 131 52
rect 123 45 126 47
rect 128 45 131 47
rect 123 43 131 45
rect 133 63 141 70
rect 133 61 136 63
rect 138 61 141 63
rect 133 43 141 61
rect 143 68 150 70
rect 143 66 146 68
rect 148 66 150 68
rect 143 60 150 66
rect 161 64 166 71
rect 143 58 146 60
rect 148 58 150 60
rect 159 62 166 64
rect 159 60 161 62
rect 163 60 166 62
rect 159 58 166 60
rect 143 43 150 58
rect 161 43 166 58
rect 168 54 176 71
rect 168 52 171 54
rect 173 52 176 54
rect 168 43 176 52
rect 178 54 186 71
rect 178 52 181 54
rect 183 52 186 54
rect 178 47 186 52
rect 178 45 181 47
rect 183 45 186 47
rect 178 43 186 45
rect 188 69 196 71
rect 188 67 191 69
rect 193 67 196 69
rect 188 57 196 67
rect 198 62 206 71
rect 198 60 201 62
rect 203 60 206 62
rect 198 57 206 60
rect 208 69 215 71
rect 208 67 211 69
rect 213 67 215 69
rect 208 62 215 67
rect 221 64 226 71
rect 208 60 211 62
rect 213 60 215 62
rect 208 57 215 60
rect 219 62 226 64
rect 219 60 221 62
rect 223 60 226 62
rect 219 58 226 60
rect 188 43 194 57
rect 221 43 226 58
rect 228 54 236 71
rect 228 52 231 54
rect 233 52 236 54
rect 228 43 236 52
rect 238 54 246 71
rect 238 52 241 54
rect 243 52 246 54
rect 238 47 246 52
rect 238 45 241 47
rect 243 45 246 47
rect 238 43 246 45
rect 248 69 255 71
rect 248 67 251 69
rect 253 67 255 69
rect 248 64 255 67
rect 248 50 257 64
rect 259 54 267 64
rect 259 52 262 54
rect 264 52 267 54
rect 259 50 267 52
rect 269 62 277 64
rect 269 60 272 62
rect 274 60 277 62
rect 319 64 324 70
rect 301 62 308 64
rect 301 61 303 62
rect 269 50 277 60
rect 292 56 297 61
rect 290 54 297 56
rect 290 52 292 54
rect 294 52 297 54
rect 248 43 255 50
rect 290 47 297 52
rect 290 45 292 47
rect 294 45 297 47
rect 290 43 297 45
rect 299 60 303 61
rect 305 60 308 62
rect 299 43 308 60
rect 317 62 324 64
rect 317 60 319 62
rect 321 60 324 62
rect 317 55 324 60
rect 317 53 319 55
rect 321 53 324 55
rect 317 51 324 53
rect 319 43 324 51
rect 326 68 334 70
rect 326 66 329 68
rect 331 66 334 68
rect 326 61 334 66
rect 326 59 329 61
rect 331 59 334 61
rect 326 43 334 59
rect 336 43 341 70
rect 343 54 351 70
rect 343 52 346 54
rect 348 52 351 54
rect 343 47 351 52
rect 343 45 346 47
rect 348 45 351 47
rect 343 43 351 45
rect 353 63 361 70
rect 353 61 356 63
rect 358 61 361 63
rect 353 43 361 61
rect 363 68 370 70
rect 363 66 366 68
rect 368 66 370 68
rect 363 60 370 66
rect 381 64 386 71
rect 363 58 366 60
rect 368 58 370 60
rect 379 62 386 64
rect 379 60 381 62
rect 383 60 386 62
rect 379 58 386 60
rect 363 43 370 58
rect 381 43 386 58
rect 388 54 396 71
rect 388 52 391 54
rect 393 52 396 54
rect 388 43 396 52
rect 398 54 406 71
rect 398 52 401 54
rect 403 52 406 54
rect 398 47 406 52
rect 398 45 401 47
rect 403 45 406 47
rect 398 43 406 45
rect 408 69 416 71
rect 408 67 411 69
rect 413 67 416 69
rect 408 57 416 67
rect 418 62 426 71
rect 418 60 421 62
rect 423 60 426 62
rect 418 57 426 60
rect 428 69 435 71
rect 428 67 431 69
rect 433 67 435 69
rect 428 62 435 67
rect 441 64 446 71
rect 428 60 431 62
rect 433 60 435 62
rect 428 57 435 60
rect 439 62 446 64
rect 439 60 441 62
rect 443 60 446 62
rect 439 58 446 60
rect 408 43 414 57
rect 441 43 446 58
rect 448 54 456 71
rect 448 52 451 54
rect 453 52 456 54
rect 448 43 456 52
rect 458 54 466 71
rect 458 52 461 54
rect 463 52 466 54
rect 458 47 466 52
rect 458 45 461 47
rect 463 45 466 47
rect 458 43 466 45
rect 468 69 475 71
rect 468 67 471 69
rect 473 67 475 69
rect 468 64 475 67
rect 468 50 477 64
rect 479 54 487 64
rect 479 52 482 54
rect 484 52 487 54
rect 479 50 487 52
rect 489 62 497 64
rect 489 60 492 62
rect 494 60 497 62
rect 489 50 497 60
rect 514 56 519 71
rect 512 54 519 56
rect 512 52 514 54
rect 516 52 519 54
rect 468 43 475 50
rect 512 47 519 52
rect 512 45 514 47
rect 516 45 519 47
rect 512 43 519 45
rect 521 69 529 71
rect 521 67 524 69
rect 526 67 529 69
rect 521 62 529 67
rect 521 60 524 62
rect 526 60 529 62
rect 521 43 529 60
rect 531 61 539 71
rect 531 59 534 61
rect 536 59 539 61
rect 531 54 539 59
rect 531 52 534 54
rect 536 52 539 54
rect 531 43 539 52
rect 541 69 555 71
rect 541 67 546 69
rect 548 68 555 69
rect 578 69 587 71
rect 548 67 557 68
rect 541 62 557 67
rect 541 60 546 62
rect 548 60 557 62
rect 541 43 557 60
rect 559 43 564 68
rect 566 59 571 68
rect 578 67 581 69
rect 583 67 587 69
rect 578 59 587 67
rect 566 50 574 59
rect 566 48 569 50
rect 571 48 574 50
rect 566 46 574 48
rect 576 46 587 59
rect 589 59 594 71
rect 589 57 596 59
rect 589 55 592 57
rect 594 55 596 57
rect 589 50 596 55
rect 589 48 592 50
rect 594 48 596 50
rect 589 46 596 48
rect 566 43 571 46
rect -210 -35 -203 -33
rect -210 -37 -208 -35
rect -206 -37 -203 -35
rect -210 -42 -203 -37
rect -210 -44 -208 -42
rect -206 -44 -203 -42
rect -210 -46 -203 -44
rect -208 -51 -203 -46
rect -201 -50 -192 -33
rect -181 -41 -176 -33
rect -201 -51 -197 -50
rect -199 -52 -197 -51
rect -195 -52 -192 -50
rect -199 -54 -192 -52
rect -183 -43 -176 -41
rect -183 -45 -181 -43
rect -179 -45 -176 -43
rect -183 -50 -176 -45
rect -183 -52 -181 -50
rect -179 -52 -176 -50
rect -183 -54 -176 -52
rect -181 -60 -176 -54
rect -174 -49 -166 -33
rect -174 -51 -171 -49
rect -169 -51 -166 -49
rect -174 -56 -166 -51
rect -174 -58 -171 -56
rect -169 -58 -166 -56
rect -174 -60 -166 -58
rect -164 -60 -159 -33
rect -157 -35 -149 -33
rect -157 -37 -154 -35
rect -152 -37 -149 -35
rect -157 -42 -149 -37
rect -157 -44 -154 -42
rect -152 -44 -149 -42
rect -157 -60 -149 -44
rect -147 -51 -139 -33
rect -147 -53 -144 -51
rect -142 -53 -139 -51
rect -147 -60 -139 -53
rect -137 -48 -130 -33
rect -119 -48 -114 -33
rect -137 -50 -134 -48
rect -132 -50 -130 -48
rect -137 -56 -130 -50
rect -121 -50 -114 -48
rect -121 -52 -119 -50
rect -117 -52 -114 -50
rect -121 -54 -114 -52
rect -137 -58 -134 -56
rect -132 -58 -130 -56
rect -137 -60 -130 -58
rect -119 -61 -114 -54
rect -112 -42 -104 -33
rect -112 -44 -109 -42
rect -107 -44 -104 -42
rect -112 -61 -104 -44
rect -102 -35 -94 -33
rect -102 -37 -99 -35
rect -97 -37 -94 -35
rect -102 -42 -94 -37
rect -102 -44 -99 -42
rect -97 -44 -94 -42
rect -102 -61 -94 -44
rect -92 -47 -86 -33
rect -92 -57 -84 -47
rect -92 -59 -89 -57
rect -87 -59 -84 -57
rect -92 -61 -84 -59
rect -82 -50 -74 -47
rect -82 -52 -79 -50
rect -77 -52 -74 -50
rect -82 -61 -74 -52
rect -72 -50 -65 -47
rect -59 -48 -54 -33
rect -72 -52 -69 -50
rect -67 -52 -65 -50
rect -72 -57 -65 -52
rect -61 -50 -54 -48
rect -61 -52 -59 -50
rect -57 -52 -54 -50
rect -61 -54 -54 -52
rect -72 -59 -69 -57
rect -67 -59 -65 -57
rect -72 -61 -65 -59
rect -59 -61 -54 -54
rect -52 -42 -44 -33
rect -52 -44 -49 -42
rect -47 -44 -44 -42
rect -52 -61 -44 -44
rect -42 -35 -34 -33
rect -42 -37 -39 -35
rect -37 -37 -34 -35
rect -42 -42 -34 -37
rect -42 -44 -39 -42
rect -37 -44 -34 -42
rect -42 -61 -34 -44
rect -32 -40 -25 -33
rect 10 -35 17 -33
rect 10 -37 12 -35
rect 14 -37 17 -35
rect -32 -54 -23 -40
rect -21 -42 -13 -40
rect -21 -44 -18 -42
rect -16 -44 -13 -42
rect -21 -54 -13 -44
rect -11 -50 -3 -40
rect 10 -42 17 -37
rect 10 -44 12 -42
rect 14 -44 17 -42
rect 10 -46 17 -44
rect -11 -52 -8 -50
rect -6 -52 -3 -50
rect 12 -51 17 -46
rect 19 -50 28 -33
rect 39 -41 44 -33
rect 19 -51 23 -50
rect -11 -54 -3 -52
rect -32 -57 -25 -54
rect -32 -59 -29 -57
rect -27 -59 -25 -57
rect 21 -52 23 -51
rect 25 -52 28 -50
rect 21 -54 28 -52
rect 37 -43 44 -41
rect 37 -45 39 -43
rect 41 -45 44 -43
rect 37 -50 44 -45
rect 37 -52 39 -50
rect 41 -52 44 -50
rect 37 -54 44 -52
rect -32 -61 -25 -59
rect 39 -60 44 -54
rect 46 -49 54 -33
rect 46 -51 49 -49
rect 51 -51 54 -49
rect 46 -56 54 -51
rect 46 -58 49 -56
rect 51 -58 54 -56
rect 46 -60 54 -58
rect 56 -60 61 -33
rect 63 -35 71 -33
rect 63 -37 66 -35
rect 68 -37 71 -35
rect 63 -42 71 -37
rect 63 -44 66 -42
rect 68 -44 71 -42
rect 63 -60 71 -44
rect 73 -51 81 -33
rect 73 -53 76 -51
rect 78 -53 81 -51
rect 73 -60 81 -53
rect 83 -48 90 -33
rect 101 -48 106 -33
rect 83 -50 86 -48
rect 88 -50 90 -48
rect 83 -56 90 -50
rect 99 -50 106 -48
rect 99 -52 101 -50
rect 103 -52 106 -50
rect 99 -54 106 -52
rect 83 -58 86 -56
rect 88 -58 90 -56
rect 83 -60 90 -58
rect 101 -61 106 -54
rect 108 -42 116 -33
rect 108 -44 111 -42
rect 113 -44 116 -42
rect 108 -61 116 -44
rect 118 -35 126 -33
rect 118 -37 121 -35
rect 123 -37 126 -35
rect 118 -42 126 -37
rect 118 -44 121 -42
rect 123 -44 126 -42
rect 118 -61 126 -44
rect 128 -47 134 -33
rect 128 -57 136 -47
rect 128 -59 131 -57
rect 133 -59 136 -57
rect 128 -61 136 -59
rect 138 -50 146 -47
rect 138 -52 141 -50
rect 143 -52 146 -50
rect 138 -61 146 -52
rect 148 -50 155 -47
rect 161 -48 166 -33
rect 148 -52 151 -50
rect 153 -52 155 -50
rect 148 -57 155 -52
rect 159 -50 166 -48
rect 159 -52 161 -50
rect 163 -52 166 -50
rect 159 -54 166 -52
rect 148 -59 151 -57
rect 153 -59 155 -57
rect 148 -61 155 -59
rect 161 -61 166 -54
rect 168 -42 176 -33
rect 168 -44 171 -42
rect 173 -44 176 -42
rect 168 -61 176 -44
rect 178 -35 186 -33
rect 178 -37 181 -35
rect 183 -37 186 -35
rect 178 -42 186 -37
rect 178 -44 181 -42
rect 183 -44 186 -42
rect 178 -61 186 -44
rect 188 -40 195 -33
rect 227 -35 234 -33
rect 227 -37 229 -35
rect 231 -37 234 -35
rect 188 -54 197 -40
rect 199 -42 207 -40
rect 199 -44 202 -42
rect 204 -44 207 -42
rect 199 -54 207 -44
rect 209 -50 217 -40
rect 227 -42 234 -37
rect 227 -44 229 -42
rect 231 -44 234 -42
rect 227 -46 234 -44
rect 209 -52 212 -50
rect 214 -52 217 -50
rect 229 -51 234 -46
rect 236 -50 245 -33
rect 256 -41 261 -33
rect 236 -51 240 -50
rect 209 -54 217 -52
rect 188 -57 195 -54
rect 188 -59 191 -57
rect 193 -59 195 -57
rect 238 -52 240 -51
rect 242 -52 245 -50
rect 238 -54 245 -52
rect 254 -43 261 -41
rect 254 -45 256 -43
rect 258 -45 261 -43
rect 254 -50 261 -45
rect 254 -52 256 -50
rect 258 -52 261 -50
rect 254 -54 261 -52
rect 188 -61 195 -59
rect 256 -60 261 -54
rect 263 -49 271 -33
rect 263 -51 266 -49
rect 268 -51 271 -49
rect 263 -56 271 -51
rect 263 -58 266 -56
rect 268 -58 271 -56
rect 263 -60 271 -58
rect 273 -60 278 -33
rect 280 -35 288 -33
rect 280 -37 283 -35
rect 285 -37 288 -35
rect 280 -42 288 -37
rect 280 -44 283 -42
rect 285 -44 288 -42
rect 280 -60 288 -44
rect 290 -51 298 -33
rect 290 -53 293 -51
rect 295 -53 298 -51
rect 290 -60 298 -53
rect 300 -48 307 -33
rect 318 -48 323 -33
rect 300 -50 303 -48
rect 305 -50 307 -48
rect 300 -56 307 -50
rect 316 -50 323 -48
rect 316 -52 318 -50
rect 320 -52 323 -50
rect 316 -54 323 -52
rect 300 -58 303 -56
rect 305 -58 307 -56
rect 300 -60 307 -58
rect 318 -61 323 -54
rect 325 -42 333 -33
rect 325 -44 328 -42
rect 330 -44 333 -42
rect 325 -61 333 -44
rect 335 -35 343 -33
rect 335 -37 338 -35
rect 340 -37 343 -35
rect 335 -42 343 -37
rect 335 -44 338 -42
rect 340 -44 343 -42
rect 335 -61 343 -44
rect 345 -47 351 -33
rect 345 -57 353 -47
rect 345 -59 348 -57
rect 350 -59 353 -57
rect 345 -61 353 -59
rect 355 -50 363 -47
rect 355 -52 358 -50
rect 360 -52 363 -50
rect 355 -61 363 -52
rect 365 -50 372 -47
rect 378 -48 383 -33
rect 365 -52 368 -50
rect 370 -52 372 -50
rect 365 -57 372 -52
rect 376 -50 383 -48
rect 376 -52 378 -50
rect 380 -52 383 -50
rect 376 -54 383 -52
rect 365 -59 368 -57
rect 370 -59 372 -57
rect 365 -61 372 -59
rect 378 -61 383 -54
rect 385 -42 393 -33
rect 385 -44 388 -42
rect 390 -44 393 -42
rect 385 -61 393 -44
rect 395 -35 403 -33
rect 395 -37 398 -35
rect 400 -37 403 -35
rect 395 -42 403 -37
rect 395 -44 398 -42
rect 400 -44 403 -42
rect 395 -61 403 -44
rect 405 -40 412 -33
rect 455 -35 462 -33
rect 455 -37 457 -35
rect 459 -37 462 -35
rect 405 -54 414 -40
rect 416 -42 424 -40
rect 416 -44 419 -42
rect 421 -44 424 -42
rect 416 -54 424 -44
rect 426 -50 434 -40
rect 455 -42 462 -37
rect 455 -44 457 -42
rect 459 -44 462 -42
rect 455 -46 462 -44
rect 426 -52 429 -50
rect 431 -52 434 -50
rect 426 -54 434 -52
rect 405 -57 412 -54
rect 405 -59 408 -57
rect 410 -59 412 -57
rect 405 -61 412 -59
rect 457 -61 462 -46
rect 464 -50 472 -33
rect 464 -52 467 -50
rect 469 -52 472 -50
rect 464 -57 472 -52
rect 464 -59 467 -57
rect 469 -59 472 -57
rect 464 -61 472 -59
rect 474 -42 482 -33
rect 474 -44 477 -42
rect 479 -44 482 -42
rect 474 -49 482 -44
rect 474 -51 477 -49
rect 479 -51 482 -49
rect 474 -61 482 -51
rect 484 -50 500 -33
rect 484 -52 489 -50
rect 491 -52 500 -50
rect 484 -57 500 -52
rect 484 -59 489 -57
rect 491 -58 500 -57
rect 502 -58 507 -33
rect 509 -36 514 -33
rect 509 -38 517 -36
rect 509 -40 512 -38
rect 514 -40 517 -38
rect 509 -49 517 -40
rect 519 -49 530 -36
rect 509 -58 514 -49
rect 521 -57 530 -49
rect 491 -59 498 -58
rect 484 -61 498 -59
rect 521 -59 524 -57
rect 526 -59 530 -57
rect 521 -61 530 -59
rect 532 -38 539 -36
rect 532 -40 535 -38
rect 537 -40 539 -38
rect 532 -45 539 -40
rect 532 -47 535 -45
rect 537 -47 539 -45
rect 532 -49 539 -47
rect 532 -61 537 -49
<< alu1 >>
rect 38 215 677 220
rect 38 213 45 215
rect 47 213 85 215
rect 87 213 128 215
rect 130 213 232 215
rect 234 213 274 215
rect 276 213 318 215
rect 320 213 387 215
rect 389 213 431 215
rect 433 213 473 215
rect 475 213 514 215
rect 516 213 557 215
rect 559 213 597 215
rect 599 213 640 215
rect 642 213 677 215
rect 38 212 677 213
rect 42 198 47 200
rect 42 196 44 198
rect 46 196 47 198
rect 42 191 47 196
rect 42 189 44 191
rect 46 189 47 191
rect 42 187 47 189
rect 74 198 78 199
rect 74 196 75 198
rect 77 196 78 198
rect 42 167 46 187
rect 74 190 78 196
rect 65 189 78 190
rect 65 187 71 189
rect 73 187 78 189
rect 65 186 78 187
rect 82 198 87 200
rect 82 196 84 198
rect 86 196 87 198
rect 82 191 87 196
rect 82 189 84 191
rect 86 189 87 191
rect 82 187 87 189
rect 114 198 118 199
rect 114 196 115 198
rect 117 196 118 198
rect 57 181 71 182
rect 57 179 61 181
rect 63 180 71 181
rect 63 179 67 180
rect 57 178 67 179
rect 69 178 71 180
rect 42 165 44 167
rect 46 165 54 167
rect 42 164 54 165
rect 42 162 48 164
rect 50 162 54 164
rect 66 169 71 178
rect 82 167 86 187
rect 114 190 118 196
rect 105 189 118 190
rect 105 187 111 189
rect 113 187 118 189
rect 105 186 118 187
rect 125 198 130 200
rect 125 196 127 198
rect 129 196 130 198
rect 125 191 130 196
rect 125 189 127 191
rect 129 189 130 191
rect 125 187 130 189
rect 157 193 161 199
rect 97 181 111 182
rect 97 179 101 181
rect 103 179 107 181
rect 109 179 111 181
rect 97 178 111 179
rect 82 165 84 167
rect 86 165 94 167
rect 82 164 94 165
rect 82 162 84 164
rect 86 162 94 164
rect 106 169 111 178
rect 125 167 129 187
rect 157 191 158 193
rect 160 191 161 193
rect 157 190 161 191
rect 148 189 161 190
rect 148 187 154 189
rect 156 187 161 189
rect 148 186 161 187
rect 229 198 234 200
rect 229 196 231 198
rect 233 196 234 198
rect 229 191 234 196
rect 229 189 231 191
rect 233 189 234 191
rect 229 187 234 189
rect 261 193 265 199
rect 140 181 154 182
rect 140 179 144 181
rect 146 179 154 181
rect 140 178 154 179
rect 125 165 127 167
rect 129 165 137 167
rect 125 164 137 165
rect 125 162 127 164
rect 129 162 137 164
rect 149 172 154 178
rect 149 170 151 172
rect 153 170 154 172
rect 149 169 154 170
rect 229 167 233 187
rect 261 191 262 193
rect 264 191 265 193
rect 261 190 265 191
rect 252 189 265 190
rect 252 187 258 189
rect 260 187 265 189
rect 252 186 265 187
rect 271 198 276 200
rect 271 196 273 198
rect 275 196 276 198
rect 271 191 276 196
rect 271 189 273 191
rect 275 189 276 191
rect 271 187 276 189
rect 303 198 307 199
rect 303 196 304 198
rect 306 196 307 198
rect 244 181 258 182
rect 244 179 248 181
rect 250 179 258 181
rect 244 178 258 179
rect 229 165 231 167
rect 233 165 241 167
rect 229 164 241 165
rect 229 162 234 164
rect 236 162 241 164
rect 253 173 258 178
rect 253 171 254 173
rect 256 171 258 173
rect 253 169 258 171
rect 271 167 275 187
rect 303 190 307 196
rect 294 189 307 190
rect 294 187 300 189
rect 302 187 307 189
rect 294 186 307 187
rect 315 198 320 200
rect 315 196 317 198
rect 319 196 320 198
rect 315 191 320 196
rect 315 189 317 191
rect 319 189 320 191
rect 315 187 320 189
rect 347 198 351 199
rect 347 196 348 198
rect 350 196 351 198
rect 286 181 300 182
rect 286 179 290 181
rect 292 179 296 181
rect 298 179 300 181
rect 286 178 300 179
rect 271 165 273 167
rect 275 165 283 167
rect 271 164 283 165
rect 271 162 272 164
rect 274 162 283 164
rect 295 169 300 178
rect 315 173 319 187
rect 315 171 316 173
rect 318 171 319 173
rect 315 167 319 171
rect 347 190 351 196
rect 338 189 351 190
rect 338 187 344 189
rect 346 187 351 189
rect 338 186 351 187
rect 384 198 389 200
rect 384 196 386 198
rect 388 196 389 198
rect 384 191 389 196
rect 384 189 386 191
rect 388 189 389 191
rect 384 187 389 189
rect 416 198 420 199
rect 416 196 417 198
rect 419 196 420 198
rect 330 181 344 182
rect 330 179 334 181
rect 336 179 344 181
rect 330 178 344 179
rect 315 165 317 167
rect 319 165 327 167
rect 42 161 54 162
rect 82 161 94 162
rect 125 161 137 162
rect 229 161 241 162
rect 271 161 283 162
rect 315 161 327 165
rect 339 173 344 178
rect 339 171 340 173
rect 342 171 344 173
rect 339 169 344 171
rect 384 167 388 187
rect 416 190 420 196
rect 407 189 420 190
rect 407 187 413 189
rect 415 187 420 189
rect 407 186 420 187
rect 428 198 433 200
rect 428 196 430 198
rect 432 196 433 198
rect 428 191 433 196
rect 428 189 430 191
rect 432 189 433 191
rect 428 187 433 189
rect 460 198 464 199
rect 460 196 461 198
rect 463 196 464 198
rect 399 181 413 182
rect 399 179 403 181
rect 405 179 413 181
rect 399 178 413 179
rect 384 165 386 167
rect 388 165 396 167
rect 384 164 396 165
rect 384 162 388 164
rect 390 162 396 164
rect 408 173 413 178
rect 408 171 409 173
rect 411 171 413 173
rect 408 169 413 171
rect 428 167 432 187
rect 460 190 464 196
rect 451 189 464 190
rect 451 187 457 189
rect 459 187 464 189
rect 451 186 464 187
rect 470 198 475 200
rect 470 196 472 198
rect 474 196 475 198
rect 470 191 475 196
rect 470 189 472 191
rect 474 189 475 191
rect 470 187 475 189
rect 502 193 506 199
rect 443 181 457 182
rect 443 179 447 181
rect 449 179 457 181
rect 443 178 457 179
rect 428 165 430 167
rect 432 165 440 167
rect 428 163 437 165
rect 439 163 440 165
rect 384 161 396 162
rect 428 161 440 163
rect 452 173 457 178
rect 452 171 453 173
rect 455 171 457 173
rect 452 169 457 171
rect 470 167 474 187
rect 502 191 503 193
rect 505 191 506 193
rect 502 190 506 191
rect 493 189 506 190
rect 493 187 499 189
rect 501 187 506 189
rect 493 186 506 187
rect 511 198 516 200
rect 511 196 513 198
rect 515 196 516 198
rect 511 191 516 196
rect 511 189 513 191
rect 515 189 516 191
rect 511 187 516 189
rect 543 197 547 199
rect 543 195 544 197
rect 546 195 547 197
rect 485 181 499 182
rect 485 179 489 181
rect 491 179 495 181
rect 497 179 499 181
rect 485 178 499 179
rect 470 165 472 167
rect 474 165 482 167
rect 470 164 482 165
rect 470 162 471 164
rect 473 162 482 164
rect 494 169 499 178
rect 511 167 515 187
rect 543 190 547 195
rect 534 189 547 190
rect 534 187 540 189
rect 542 187 547 189
rect 534 186 547 187
rect 554 198 559 200
rect 554 196 556 198
rect 558 196 559 198
rect 554 191 559 196
rect 554 189 556 191
rect 558 189 559 191
rect 554 187 559 189
rect 586 198 590 199
rect 586 196 587 198
rect 589 196 590 198
rect 526 181 540 182
rect 526 179 530 181
rect 532 179 540 181
rect 526 178 540 179
rect 511 165 513 167
rect 515 165 523 167
rect 511 164 523 165
rect 511 162 519 164
rect 521 162 523 164
rect 535 173 540 178
rect 535 171 536 173
rect 538 171 540 173
rect 535 169 540 171
rect 554 167 558 187
rect 586 190 590 196
rect 577 189 590 190
rect 577 187 583 189
rect 585 187 590 189
rect 577 186 590 187
rect 594 198 599 200
rect 594 196 596 198
rect 598 196 599 198
rect 594 191 599 196
rect 594 189 596 191
rect 598 189 599 191
rect 594 187 599 189
rect 626 193 630 199
rect 569 181 583 182
rect 569 179 573 181
rect 575 179 579 181
rect 581 179 583 181
rect 569 178 583 179
rect 554 165 556 167
rect 558 165 566 167
rect 554 164 566 165
rect 554 162 562 164
rect 564 162 566 164
rect 578 169 583 178
rect 594 167 598 187
rect 626 191 627 193
rect 629 191 630 193
rect 626 190 630 191
rect 617 189 630 190
rect 617 187 623 189
rect 625 187 630 189
rect 617 186 630 187
rect 637 198 642 200
rect 637 196 639 198
rect 641 196 642 198
rect 637 191 642 196
rect 637 189 639 191
rect 641 189 642 191
rect 637 187 642 189
rect 669 198 673 199
rect 669 196 670 198
rect 672 196 673 198
rect 609 181 623 182
rect 609 179 613 181
rect 615 179 623 181
rect 609 178 623 179
rect 594 165 596 167
rect 598 165 606 167
rect 594 164 606 165
rect 594 162 602 164
rect 604 162 606 164
rect 618 172 623 178
rect 618 170 620 172
rect 622 170 623 172
rect 618 169 623 170
rect 637 167 641 187
rect 669 190 673 196
rect 660 189 673 190
rect 660 187 666 189
rect 668 187 673 189
rect 660 186 673 187
rect 652 181 666 182
rect 652 179 656 181
rect 658 179 666 181
rect 652 178 666 179
rect 637 165 639 167
rect 641 165 649 167
rect 470 161 482 162
rect 511 161 523 162
rect 554 161 566 162
rect 594 161 606 162
rect 637 161 649 165
rect 661 172 666 178
rect 661 170 663 172
rect 665 170 666 172
rect 661 169 666 170
rect 38 155 677 156
rect 38 153 45 155
rect 47 153 55 155
rect 57 153 85 155
rect 87 153 95 155
rect 97 153 128 155
rect 130 153 138 155
rect 140 153 232 155
rect 234 153 242 155
rect 244 153 274 155
rect 276 153 284 155
rect 286 153 318 155
rect 320 153 328 155
rect 330 153 387 155
rect 389 153 397 155
rect 399 153 431 155
rect 433 153 441 155
rect 443 153 473 155
rect 475 153 483 155
rect 485 153 514 155
rect 516 153 524 155
rect 526 153 557 155
rect 559 153 567 155
rect 569 153 597 155
rect 599 153 607 155
rect 609 153 640 155
rect 642 153 650 155
rect 652 153 677 155
rect 38 149 677 153
rect -79 148 677 149
rect -79 144 641 148
rect -79 142 -72 144
rect -70 142 -62 144
rect -60 142 -30 144
rect -28 142 -20 144
rect -18 142 109 144
rect 111 142 121 144
rect 123 142 143 144
rect 145 142 197 144
rect 199 142 259 144
rect 261 142 314 144
rect 316 142 327 144
rect 329 142 339 144
rect 341 142 361 144
rect 363 142 415 144
rect 417 142 477 144
rect 479 142 532 144
rect 534 142 641 144
rect -79 141 641 142
rect -75 132 -63 136
rect -75 130 -73 132
rect -71 130 -63 132
rect -33 132 -21 136
rect -75 110 -71 130
rect -33 130 -31 132
rect -29 130 -21 132
rect 14 134 36 135
rect 14 132 17 134
rect 19 132 36 134
rect 14 131 36 132
rect 94 134 99 136
rect 94 132 95 134
rect 97 132 99 134
rect -51 119 -46 128
rect -75 108 -70 110
rect -75 106 -73 108
rect -71 106 -70 108
rect -75 105 -70 106
rect -75 103 -74 105
rect -72 103 -70 105
rect -75 101 -70 103
rect -75 99 -73 101
rect -71 99 -70 101
rect -60 118 -46 119
rect -60 116 -59 118
rect -57 116 -56 118
rect -54 116 -46 118
rect -60 115 -46 116
rect -52 110 -39 111
rect -52 108 -46 110
rect -44 108 -42 110
rect -40 108 -39 110
rect -52 107 -39 108
rect -75 97 -70 99
rect -43 98 -39 107
rect -33 110 -29 130
rect -9 119 -4 128
rect -33 108 -28 110
rect -33 106 -31 108
rect -29 106 -28 108
rect -33 104 -28 106
rect -33 102 -32 104
rect -30 102 -28 104
rect -33 101 -28 102
rect -33 99 -31 101
rect -29 99 -28 101
rect -18 118 -4 119
rect -18 116 -17 118
rect -15 116 -14 118
rect -12 116 -4 118
rect -18 115 -4 116
rect 14 111 18 131
rect 47 126 51 128
rect 47 124 48 126
rect 50 124 51 126
rect -10 110 3 111
rect -10 108 -4 110
rect -2 108 0 110
rect 2 108 3 110
rect -10 107 3 108
rect -33 97 -28 99
rect -1 98 3 107
rect 14 109 20 111
rect 14 107 17 109
rect 19 107 20 109
rect 14 105 20 107
rect 14 103 16 105
rect 18 103 20 105
rect 14 102 20 103
rect 14 100 17 102
rect 19 100 20 102
rect 14 98 20 100
rect 47 119 51 124
rect 94 130 99 132
rect 63 119 71 120
rect 38 118 53 119
rect 38 116 42 118
rect 44 116 49 118
rect 51 116 53 118
rect 38 115 53 116
rect 63 117 64 119
rect 66 118 71 119
rect 66 117 68 118
rect 63 116 68 117
rect 70 116 71 118
rect 63 114 71 116
rect 63 111 68 114
rect 30 107 68 111
rect 95 108 99 130
rect 94 106 99 108
rect 94 104 95 106
rect 97 104 99 106
rect 94 99 99 104
rect 94 97 95 99
rect 97 97 99 99
rect 106 127 110 136
rect 195 134 219 135
rect 195 132 215 134
rect 217 132 219 134
rect 195 131 219 132
rect 106 125 108 127
rect 106 109 110 125
rect 114 127 118 128
rect 114 125 115 127
rect 117 125 118 127
rect 146 127 165 128
rect 146 126 161 127
rect 114 120 118 125
rect 146 124 147 126
rect 149 125 161 126
rect 163 125 165 127
rect 149 124 165 125
rect 146 123 165 124
rect 169 126 183 127
rect 169 124 180 126
rect 182 124 183 126
rect 169 123 183 124
rect 114 118 126 120
rect 114 116 115 118
rect 117 116 126 118
rect 114 114 126 116
rect 130 118 142 120
rect 130 116 139 118
rect 141 116 142 118
rect 130 114 142 116
rect 106 107 108 109
rect 106 104 110 107
rect 130 106 134 114
rect 146 111 150 123
rect 169 119 173 123
rect 161 118 173 119
rect 161 116 165 118
rect 167 116 173 118
rect 161 115 173 116
rect 177 118 183 119
rect 177 116 179 118
rect 181 116 183 118
rect 177 111 183 116
rect 146 109 166 111
rect 146 107 162 109
rect 164 107 166 109
rect 106 102 118 104
rect 106 100 108 102
rect 110 100 115 102
rect 117 100 118 102
rect 106 98 118 100
rect 94 95 99 97
rect 86 94 99 95
rect 86 92 87 94
rect 89 92 99 94
rect 86 91 99 92
rect 161 102 166 107
rect 161 100 162 102
rect 164 100 166 102
rect 161 98 166 100
rect 170 106 183 111
rect 170 101 174 106
rect 170 99 171 101
rect 173 99 174 101
rect 195 103 199 131
rect 243 124 247 126
rect 243 122 244 124
rect 246 122 247 124
rect 243 121 247 122
rect 243 119 244 121
rect 246 119 247 121
rect 195 102 211 103
rect 195 100 200 102
rect 202 100 207 102
rect 209 100 211 102
rect 195 99 211 100
rect 170 98 174 99
rect 243 105 247 119
rect 234 104 247 105
rect 234 102 240 104
rect 242 102 247 104
rect 234 99 247 102
rect 298 120 304 127
rect 291 119 304 120
rect 291 117 292 119
rect 294 117 304 119
rect 291 114 304 117
rect 324 127 328 136
rect 413 134 437 135
rect 413 132 433 134
rect 435 132 437 134
rect 413 131 437 132
rect 324 125 326 127
rect 315 119 319 120
rect 315 117 316 119
rect 318 117 319 119
rect 315 113 319 117
rect 314 111 319 113
rect 314 109 315 111
rect 317 109 319 111
rect 314 107 319 109
rect 315 103 319 107
rect 306 102 319 103
rect 306 100 308 102
rect 310 100 319 102
rect 306 98 319 100
rect 324 109 328 125
rect 332 127 336 128
rect 332 125 333 127
rect 335 125 336 127
rect 364 127 383 128
rect 364 126 379 127
rect 332 120 336 125
rect 364 124 365 126
rect 367 125 379 126
rect 381 125 383 127
rect 367 124 383 125
rect 364 123 383 124
rect 387 126 401 127
rect 387 124 388 126
rect 390 124 398 126
rect 400 124 401 126
rect 387 123 401 124
rect 332 118 344 120
rect 332 116 333 118
rect 335 116 344 118
rect 332 114 344 116
rect 348 118 360 120
rect 348 116 357 118
rect 359 116 360 118
rect 348 114 360 116
rect 324 107 326 109
rect 324 104 328 107
rect 348 106 352 114
rect 364 111 368 123
rect 387 119 391 123
rect 379 118 391 119
rect 379 116 383 118
rect 385 116 391 118
rect 379 115 391 116
rect 395 118 401 119
rect 395 116 397 118
rect 399 116 401 118
rect 395 111 401 116
rect 364 109 384 111
rect 364 107 380 109
rect 382 107 384 109
rect 324 102 336 104
rect 324 100 326 102
rect 328 100 333 102
rect 335 100 336 102
rect 324 98 336 100
rect 379 102 384 107
rect 379 100 380 102
rect 382 100 384 102
rect 379 98 384 100
rect 388 106 401 111
rect 388 101 392 106
rect 388 99 389 101
rect 391 99 392 101
rect 413 103 417 131
rect 552 134 574 135
rect 552 132 555 134
rect 557 132 574 134
rect 552 131 574 132
rect 632 134 637 136
rect 632 132 633 134
rect 635 132 637 134
rect 461 124 465 126
rect 461 122 462 124
rect 464 122 465 124
rect 461 121 465 122
rect 461 119 462 121
rect 464 119 465 121
rect 413 102 429 103
rect 413 100 421 102
rect 423 100 425 102
rect 427 100 429 102
rect 413 99 429 100
rect 388 98 392 99
rect 461 105 465 119
rect 452 104 465 105
rect 452 102 458 104
rect 460 102 465 104
rect 452 99 465 102
rect 516 120 522 127
rect 509 119 522 120
rect 509 117 510 119
rect 512 117 522 119
rect 509 114 522 117
rect 533 119 537 120
rect 533 117 534 119
rect 536 117 537 119
rect 533 113 537 117
rect 532 111 537 113
rect 532 109 533 111
rect 535 109 537 111
rect 532 107 537 109
rect 533 103 537 107
rect 524 102 537 103
rect 524 100 526 102
rect 528 100 537 102
rect 524 98 537 100
rect 552 111 556 131
rect 585 126 589 128
rect 585 124 586 126
rect 588 124 589 126
rect 552 109 558 111
rect 552 107 555 109
rect 557 107 558 109
rect 552 106 558 107
rect 552 104 554 106
rect 556 104 558 106
rect 552 102 558 104
rect 552 100 555 102
rect 557 100 558 102
rect 552 98 558 100
rect 585 119 589 124
rect 632 130 637 132
rect 601 119 609 120
rect 576 118 591 119
rect 576 116 580 118
rect 582 116 587 118
rect 589 116 591 118
rect 576 115 591 116
rect 601 117 602 119
rect 604 118 609 119
rect 604 117 606 118
rect 601 116 606 117
rect 608 116 609 118
rect 601 114 609 116
rect 601 111 606 114
rect 568 107 606 111
rect 633 108 637 130
rect 632 106 637 108
rect 632 104 633 106
rect 635 104 637 106
rect 632 99 637 104
rect 632 97 633 99
rect 635 97 637 99
rect 632 95 637 97
rect 624 91 637 95
rect -79 84 641 85
rect -79 82 -72 84
rect -70 82 -30 84
rect -28 82 109 84
rect 111 82 121 84
rect 123 82 314 84
rect 316 82 327 84
rect 329 82 339 84
rect 341 82 532 84
rect 534 82 641 84
rect -79 77 641 82
rect -196 72 600 77
rect -196 70 -189 72
rect -187 70 -145 72
rect -143 70 -133 72
rect -131 70 60 72
rect 62 70 73 72
rect 75 70 85 72
rect 87 70 278 72
rect 280 70 293 72
rect 295 70 305 72
rect 307 70 498 72
rect 500 70 600 72
rect -196 69 600 70
rect -192 55 -187 57
rect -192 53 -190 55
rect -188 53 -187 55
rect -192 48 -187 53
rect -192 46 -190 48
rect -188 46 -187 48
rect -192 44 -187 46
rect -160 55 -156 56
rect -160 53 -159 55
rect -157 53 -156 55
rect -192 24 -188 44
rect -160 47 -156 53
rect -169 46 -156 47
rect -169 44 -163 46
rect -161 44 -156 46
rect -169 43 -156 44
rect -148 54 -136 56
rect -148 52 -146 54
rect -144 52 -136 54
rect -148 50 -136 52
rect -93 54 -88 56
rect -93 52 -92 54
rect -90 52 -88 54
rect -148 47 -144 50
rect -148 45 -146 47
rect -177 38 -163 39
rect -177 36 -176 38
rect -174 36 -173 38
rect -171 36 -163 38
rect -177 35 -163 36
rect -192 22 -190 24
rect -188 22 -180 24
rect -192 21 -180 22
rect -192 19 -191 21
rect -189 19 -180 21
rect -168 26 -163 35
rect -148 29 -144 45
rect -124 40 -120 48
rect -93 47 -88 52
rect -108 45 -92 47
rect -90 45 -88 47
rect -108 43 -88 45
rect -84 55 -80 56
rect -84 53 -83 55
rect -81 53 -80 55
rect -84 48 -80 53
rect -59 54 -43 55
rect -59 52 -47 54
rect -45 52 -43 54
rect -59 51 -43 52
rect -84 43 -71 48
rect -140 38 -128 40
rect -140 36 -139 38
rect -137 36 -128 38
rect -140 34 -128 36
rect -124 38 -112 40
rect -124 36 -115 38
rect -113 36 -112 38
rect -124 34 -112 36
rect -148 27 -146 29
rect -148 21 -144 27
rect -140 29 -136 34
rect -140 27 -139 29
rect -137 27 -136 29
rect -108 31 -104 43
rect -93 38 -81 39
rect -93 36 -89 38
rect -87 36 -81 38
rect -93 35 -81 36
rect -77 38 -71 43
rect -77 36 -75 38
rect -73 36 -71 38
rect -77 35 -71 36
rect -85 31 -81 35
rect -108 30 -89 31
rect -108 28 -107 30
rect -105 29 -89 30
rect -105 28 -93 29
rect -140 26 -136 27
rect -108 27 -93 28
rect -91 27 -89 29
rect -85 30 -71 31
rect -85 28 -74 30
rect -72 28 -71 30
rect -85 27 -71 28
rect -108 26 -89 27
rect -148 19 -147 21
rect -145 19 -144 21
rect -192 18 -180 19
rect -148 18 -144 19
rect -59 23 -55 51
rect -20 52 -7 55
rect -20 50 -14 52
rect -12 50 -7 52
rect -20 49 -7 50
rect -59 22 -35 23
rect -59 20 -47 22
rect -45 20 -39 22
rect -37 20 -35 22
rect -59 19 -35 20
rect -11 35 -7 49
rect -11 33 -10 35
rect -8 33 -7 35
rect -11 32 -7 33
rect -11 30 -10 32
rect -8 30 -7 32
rect -11 28 -7 30
rect 52 54 65 56
rect 52 52 54 54
rect 56 52 65 54
rect 52 51 65 52
rect 61 47 65 51
rect 37 37 50 40
rect 37 35 38 37
rect 40 35 50 37
rect 37 34 50 35
rect 44 27 50 34
rect 60 45 65 47
rect 60 43 61 45
rect 63 43 65 45
rect 60 41 65 43
rect 61 34 65 41
rect 70 54 82 56
rect 70 52 72 54
rect 74 52 82 54
rect 70 50 82 52
rect 125 54 130 56
rect 125 52 126 54
rect 128 52 130 54
rect 70 47 74 50
rect 70 45 72 47
rect 70 29 74 45
rect 94 40 98 48
rect 125 47 130 52
rect 110 45 126 47
rect 128 45 130 47
rect 110 43 130 45
rect 134 55 138 56
rect 134 53 135 55
rect 137 53 138 55
rect 134 48 138 53
rect 159 54 175 55
rect 159 52 171 54
rect 173 52 175 54
rect 159 51 175 52
rect 134 43 147 48
rect 78 38 90 40
rect 78 36 79 38
rect 81 36 90 38
rect 78 34 90 36
rect 94 38 106 40
rect 94 36 103 38
rect 105 36 106 38
rect 94 34 106 36
rect 70 27 72 29
rect 70 21 74 27
rect 78 29 82 34
rect 78 27 79 29
rect 81 27 82 29
rect 110 31 114 43
rect 125 38 137 39
rect 125 36 129 38
rect 131 36 137 38
rect 125 35 137 36
rect 141 38 147 43
rect 141 36 143 38
rect 145 36 147 38
rect 141 35 147 36
rect 133 31 137 35
rect 110 30 129 31
rect 110 28 111 30
rect 113 29 129 30
rect 113 28 125 29
rect 78 26 82 27
rect 110 27 125 28
rect 127 27 129 29
rect 133 30 147 31
rect 133 28 144 30
rect 146 28 147 30
rect 133 27 147 28
rect 110 26 129 27
rect 70 19 71 21
rect 73 19 74 21
rect 70 18 74 19
rect 159 23 163 51
rect 198 52 211 55
rect 198 50 204 52
rect 206 50 211 52
rect 198 49 211 50
rect 159 22 183 23
rect 159 20 170 22
rect 172 20 179 22
rect 181 20 183 22
rect 159 19 183 20
rect 207 35 211 49
rect 207 33 208 35
rect 210 33 211 35
rect 207 32 211 33
rect 207 30 208 32
rect 210 30 211 32
rect 207 28 211 30
rect 270 54 283 56
rect 270 52 272 54
rect 274 52 283 54
rect 270 51 283 52
rect 279 47 283 51
rect 255 37 268 40
rect 255 35 256 37
rect 258 35 268 37
rect 255 34 268 35
rect 262 27 268 34
rect 278 45 283 47
rect 278 43 279 45
rect 281 43 283 45
rect 278 41 283 43
rect 279 34 283 41
rect 290 54 302 56
rect 290 52 292 54
rect 294 52 302 54
rect 290 50 302 52
rect 583 59 596 63
rect 345 54 350 56
rect 345 52 346 54
rect 348 52 350 54
rect 290 47 294 50
rect 290 45 292 47
rect 290 29 294 45
rect 314 40 318 48
rect 345 47 350 52
rect 330 45 346 47
rect 348 45 350 47
rect 330 43 350 45
rect 354 55 358 56
rect 354 53 355 55
rect 357 53 358 55
rect 354 48 358 53
rect 379 54 395 55
rect 379 52 391 54
rect 393 52 395 54
rect 379 51 395 52
rect 354 43 367 48
rect 298 38 310 40
rect 298 36 299 38
rect 301 36 310 38
rect 298 34 310 36
rect 314 38 326 40
rect 314 36 323 38
rect 325 36 326 38
rect 314 34 326 36
rect 290 27 292 29
rect 290 21 294 27
rect 298 29 302 34
rect 298 27 299 29
rect 301 27 302 29
rect 330 31 334 43
rect 345 38 357 39
rect 345 36 346 38
rect 348 36 349 38
rect 351 36 357 38
rect 345 35 357 36
rect 361 38 367 43
rect 361 36 363 38
rect 365 36 367 38
rect 361 35 367 36
rect 353 31 357 35
rect 330 30 349 31
rect 330 28 331 30
rect 333 29 349 30
rect 333 28 345 29
rect 298 26 302 27
rect 330 27 345 28
rect 347 27 349 29
rect 353 30 367 31
rect 353 28 364 30
rect 366 28 367 30
rect 353 27 367 28
rect 330 26 349 27
rect 290 19 291 21
rect 293 19 294 21
rect 290 18 294 19
rect 379 23 383 51
rect 418 52 431 55
rect 418 50 424 52
rect 426 50 431 52
rect 418 49 431 50
rect 379 22 403 23
rect 379 20 391 22
rect 393 20 399 22
rect 401 20 403 22
rect 379 19 403 20
rect 427 35 431 49
rect 427 33 428 35
rect 430 33 431 35
rect 427 32 431 33
rect 427 30 428 32
rect 430 30 431 32
rect 427 28 431 30
rect 490 54 503 56
rect 490 52 492 54
rect 494 52 503 54
rect 490 51 503 52
rect 499 47 503 51
rect 475 37 488 40
rect 475 35 476 37
rect 478 35 488 37
rect 475 34 488 35
rect 482 27 488 34
rect 498 45 503 47
rect 498 43 499 45
rect 501 43 503 45
rect 498 41 503 43
rect 499 34 503 41
rect 511 54 517 56
rect 591 57 596 59
rect 591 55 592 57
rect 594 55 596 57
rect 511 52 514 54
rect 516 52 517 54
rect 511 47 517 52
rect 511 45 514 47
rect 516 45 517 47
rect 511 43 517 45
rect 511 25 515 43
rect 527 46 565 47
rect 527 44 553 46
rect 555 44 565 46
rect 527 43 565 44
rect 560 40 565 43
rect 535 38 550 39
rect 535 36 536 38
rect 538 36 539 38
rect 541 36 546 38
rect 548 36 550 38
rect 535 35 550 36
rect 560 38 568 40
rect 560 36 565 38
rect 567 36 568 38
rect 511 23 512 25
rect 514 23 515 25
rect 544 26 548 35
rect 560 34 568 36
rect 591 50 596 55
rect 591 48 592 50
rect 594 48 596 50
rect 591 46 596 48
rect 511 22 533 23
rect 511 20 514 22
rect 516 20 533 22
rect 511 19 533 20
rect 592 24 596 46
rect 591 22 596 24
rect 591 20 592 22
rect 594 20 596 22
rect 591 18 596 20
rect -196 12 600 13
rect -196 10 -189 12
rect -187 10 -179 12
rect -177 10 -145 12
rect -143 10 -133 12
rect -131 10 -111 12
rect -109 10 -57 12
rect -55 10 5 12
rect 7 10 60 12
rect 62 10 73 12
rect 75 10 85 12
rect 87 10 107 12
rect 109 10 161 12
rect 163 10 223 12
rect 225 10 278 12
rect 280 10 293 12
rect 295 10 305 12
rect 307 10 327 12
rect 329 10 381 12
rect 383 10 443 12
rect 445 10 498 12
rect 500 10 600 12
rect -196 5 600 10
rect -214 0 543 5
rect -214 -2 -207 0
rect -205 -2 -195 0
rect -193 -2 -173 0
rect -171 -2 -119 0
rect -117 -2 -57 0
rect -55 -2 -2 0
rect 0 -2 13 0
rect 15 -2 25 0
rect 27 -2 47 0
rect 49 -2 101 0
rect 103 -2 163 0
rect 165 -2 218 0
rect 220 -2 230 0
rect 232 -2 242 0
rect 244 -2 264 0
rect 266 -2 318 0
rect 320 -2 380 0
rect 382 -2 435 0
rect 437 -2 543 0
rect -214 -3 543 -2
rect -210 -17 -206 -8
rect -121 -10 -97 -9
rect -121 -12 -101 -10
rect -99 -12 -97 -10
rect -121 -13 -97 -12
rect -210 -19 -208 -17
rect -210 -35 -206 -19
rect -202 -17 -198 -16
rect -202 -19 -201 -17
rect -199 -19 -198 -17
rect -170 -17 -151 -16
rect -170 -18 -155 -17
rect -202 -24 -198 -19
rect -170 -20 -169 -18
rect -167 -19 -155 -18
rect -153 -19 -151 -17
rect -167 -20 -151 -19
rect -170 -21 -151 -20
rect -147 -18 -133 -17
rect -147 -20 -136 -18
rect -134 -20 -133 -18
rect -147 -21 -133 -20
rect -202 -26 -190 -24
rect -202 -28 -201 -26
rect -199 -28 -190 -26
rect -202 -30 -190 -28
rect -186 -26 -174 -24
rect -186 -28 -177 -26
rect -175 -28 -174 -26
rect -186 -30 -174 -28
rect -210 -37 -208 -35
rect -210 -40 -206 -37
rect -186 -38 -182 -30
rect -170 -33 -166 -21
rect -147 -25 -143 -21
rect -155 -26 -143 -25
rect -155 -28 -151 -26
rect -149 -28 -143 -26
rect -155 -29 -143 -28
rect -139 -26 -133 -25
rect -139 -28 -137 -26
rect -135 -28 -133 -26
rect -139 -33 -133 -28
rect -170 -35 -150 -33
rect -170 -37 -154 -35
rect -152 -37 -150 -35
rect -210 -42 -198 -40
rect -210 -44 -208 -42
rect -206 -44 -198 -42
rect -210 -46 -198 -44
rect -155 -42 -150 -37
rect -155 -44 -154 -42
rect -152 -44 -150 -42
rect -155 -46 -150 -44
rect -146 -38 -133 -33
rect -146 -43 -142 -38
rect -146 -45 -145 -43
rect -143 -45 -142 -43
rect -121 -41 -117 -13
rect -73 -20 -69 -18
rect -73 -22 -72 -20
rect -70 -22 -69 -20
rect -73 -23 -69 -22
rect -73 -25 -72 -23
rect -70 -25 -69 -23
rect -121 -42 -105 -41
rect -121 -44 -109 -42
rect -107 -44 -105 -42
rect -121 -45 -105 -44
rect -146 -46 -142 -45
rect -73 -39 -69 -25
rect -82 -40 -69 -39
rect -82 -42 -76 -40
rect -74 -42 -69 -40
rect -82 -45 -69 -42
rect -18 -24 -12 -17
rect -25 -25 -12 -24
rect -25 -27 -24 -25
rect -22 -27 -12 -25
rect -25 -30 -12 -27
rect 10 -17 14 -8
rect 99 -10 123 -9
rect 99 -12 119 -10
rect 121 -12 123 -10
rect 99 -13 123 -12
rect 10 -19 12 -17
rect -1 -31 3 -24
rect -2 -33 3 -31
rect -2 -35 -1 -33
rect 1 -35 3 -33
rect -2 -37 3 -35
rect -1 -41 3 -37
rect -10 -42 3 -41
rect -10 -44 -8 -42
rect -6 -44 3 -42
rect -10 -46 3 -44
rect 10 -35 14 -19
rect 18 -17 22 -16
rect 18 -19 19 -17
rect 21 -19 22 -17
rect 50 -17 69 -16
rect 50 -18 65 -17
rect 18 -24 22 -19
rect 50 -20 51 -18
rect 53 -19 65 -18
rect 67 -19 69 -17
rect 53 -20 69 -19
rect 50 -21 69 -20
rect 73 -18 87 -17
rect 73 -20 84 -18
rect 86 -20 87 -18
rect 73 -21 87 -20
rect 18 -26 30 -24
rect 18 -28 19 -26
rect 21 -28 30 -26
rect 18 -30 30 -28
rect 34 -26 46 -24
rect 34 -28 43 -26
rect 45 -28 46 -26
rect 34 -30 46 -28
rect 10 -37 12 -35
rect 10 -39 14 -37
rect 10 -41 11 -39
rect 13 -40 14 -39
rect 34 -38 38 -30
rect 50 -33 54 -21
rect 73 -25 77 -21
rect 65 -26 77 -25
rect 65 -28 69 -26
rect 71 -28 77 -26
rect 65 -29 77 -28
rect 81 -26 87 -25
rect 81 -28 83 -26
rect 85 -28 87 -26
rect 81 -33 87 -28
rect 50 -35 70 -33
rect 50 -37 66 -35
rect 68 -37 70 -35
rect 13 -41 22 -40
rect 10 -42 22 -41
rect 10 -44 12 -42
rect 14 -44 22 -42
rect 10 -46 22 -44
rect 65 -42 70 -37
rect 65 -44 66 -42
rect 68 -44 70 -42
rect 65 -46 70 -44
rect 74 -38 87 -33
rect 74 -43 78 -38
rect 74 -45 75 -43
rect 77 -45 78 -43
rect 99 -41 103 -13
rect 147 -20 151 -18
rect 147 -22 148 -20
rect 150 -22 151 -20
rect 147 -23 151 -22
rect 147 -25 148 -23
rect 150 -25 151 -23
rect 99 -42 115 -41
rect 99 -44 111 -42
rect 113 -44 115 -42
rect 99 -45 115 -44
rect 74 -46 78 -45
rect 147 -39 151 -25
rect 138 -40 151 -39
rect 138 -42 144 -40
rect 146 -42 151 -40
rect 138 -45 151 -42
rect 202 -24 208 -17
rect 195 -25 208 -24
rect 195 -27 196 -25
rect 198 -27 208 -25
rect 195 -30 208 -27
rect 227 -17 231 -8
rect 316 -10 340 -9
rect 316 -12 336 -10
rect 338 -12 340 -10
rect 316 -13 340 -12
rect 227 -19 229 -17
rect 219 -31 223 -24
rect 218 -33 223 -31
rect 218 -35 219 -33
rect 221 -35 223 -33
rect 218 -37 223 -35
rect 219 -41 223 -37
rect 210 -42 223 -41
rect 210 -44 212 -42
rect 214 -44 223 -42
rect 210 -46 223 -44
rect 227 -35 231 -19
rect 235 -17 239 -16
rect 235 -19 236 -17
rect 238 -19 239 -17
rect 267 -17 286 -16
rect 267 -18 282 -17
rect 235 -24 239 -19
rect 267 -20 268 -18
rect 270 -19 282 -18
rect 284 -19 286 -17
rect 270 -20 286 -19
rect 267 -21 286 -20
rect 290 -18 304 -17
rect 290 -20 291 -18
rect 293 -20 301 -18
rect 303 -20 304 -18
rect 290 -21 304 -20
rect 235 -26 247 -24
rect 235 -28 236 -26
rect 238 -28 247 -26
rect 235 -30 247 -28
rect 251 -26 263 -24
rect 251 -28 260 -26
rect 262 -28 263 -26
rect 251 -30 263 -28
rect 227 -37 229 -35
rect 227 -38 231 -37
rect 227 -40 228 -38
rect 230 -40 231 -38
rect 251 -38 255 -30
rect 267 -33 271 -21
rect 290 -25 294 -21
rect 282 -26 294 -25
rect 282 -28 286 -26
rect 288 -28 294 -26
rect 282 -29 294 -28
rect 298 -26 304 -25
rect 298 -28 300 -26
rect 302 -28 304 -26
rect 298 -33 304 -28
rect 267 -35 287 -33
rect 267 -37 283 -35
rect 285 -37 287 -35
rect 227 -42 239 -40
rect 227 -44 229 -42
rect 231 -44 239 -42
rect 227 -46 239 -44
rect 282 -42 287 -37
rect 282 -44 283 -42
rect 285 -44 287 -42
rect 282 -46 287 -44
rect 291 -38 304 -33
rect 291 -43 295 -38
rect 291 -45 292 -43
rect 294 -45 295 -43
rect 316 -41 320 -13
rect 454 -10 476 -9
rect 454 -12 457 -10
rect 459 -12 476 -10
rect 454 -13 476 -12
rect 534 -10 539 -8
rect 534 -12 535 -10
rect 537 -12 539 -10
rect 364 -20 368 -18
rect 364 -22 365 -20
rect 367 -22 368 -20
rect 364 -23 368 -22
rect 364 -25 365 -23
rect 367 -25 368 -23
rect 316 -42 332 -41
rect 316 -44 328 -42
rect 330 -44 332 -42
rect 316 -45 332 -44
rect 291 -46 295 -45
rect 364 -39 368 -25
rect 355 -40 368 -39
rect 355 -42 361 -40
rect 363 -42 368 -40
rect 355 -45 368 -42
rect 419 -24 425 -17
rect 412 -25 425 -24
rect 412 -27 413 -25
rect 415 -27 425 -25
rect 412 -30 425 -27
rect 436 -31 440 -24
rect 435 -33 440 -31
rect 435 -35 436 -33
rect 438 -35 440 -33
rect 435 -37 440 -35
rect 436 -41 440 -37
rect 427 -42 440 -41
rect 427 -44 429 -42
rect 431 -44 440 -42
rect 427 -46 440 -44
rect 454 -33 458 -13
rect 487 -17 491 -16
rect 487 -19 488 -17
rect 490 -19 491 -17
rect 454 -35 460 -33
rect 454 -37 457 -35
rect 459 -37 460 -35
rect 454 -39 460 -37
rect 454 -41 455 -39
rect 457 -41 460 -39
rect 454 -42 460 -41
rect 454 -44 457 -42
rect 459 -44 460 -42
rect 454 -46 460 -44
rect 487 -25 491 -19
rect 534 -14 539 -12
rect 478 -26 493 -25
rect 478 -28 482 -26
rect 484 -28 489 -26
rect 491 -28 493 -26
rect 478 -29 493 -28
rect 503 -26 511 -24
rect 503 -28 508 -26
rect 510 -28 511 -26
rect 503 -30 511 -28
rect 503 -33 508 -30
rect 470 -34 508 -33
rect 470 -36 472 -34
rect 474 -36 508 -34
rect 470 -37 508 -36
rect 535 -36 539 -14
rect 534 -38 539 -36
rect 534 -40 535 -38
rect 537 -40 539 -38
rect 534 -45 539 -40
rect 534 -47 535 -45
rect 537 -47 539 -45
rect 534 -49 539 -47
rect 526 -53 539 -49
rect -214 -60 543 -59
rect -214 -62 -207 -60
rect -205 -62 -195 -60
rect -193 -62 -2 -60
rect 0 -62 13 -60
rect 15 -62 25 -60
rect 27 -62 218 -60
rect 220 -62 230 -60
rect 232 -62 242 -60
rect 244 -62 435 -60
rect 437 -62 543 -60
rect -214 -67 543 -62
<< alu2 >>
rect -160 213 -156 214
rect -160 211 -159 213
rect -157 211 -156 213
rect -177 150 -173 152
rect -177 148 -176 150
rect -174 148 -173 150
rect -177 38 -173 148
rect -160 55 -156 211
rect -43 213 -39 214
rect -43 211 -42 213
rect -40 211 -39 213
rect -60 161 -56 162
rect -60 159 -59 161
rect -57 159 -56 161
rect -60 118 -56 159
rect -60 116 -59 118
rect -57 116 -56 118
rect -60 115 -56 116
rect -43 110 -39 211
rect 114 213 118 214
rect 114 211 115 213
rect 117 211 118 213
rect -1 202 3 203
rect -1 200 0 202
rect 2 200 3 202
rect -18 150 -14 152
rect -18 148 -17 150
rect -15 148 -14 150
rect -18 118 -14 148
rect -18 116 -17 118
rect -15 116 -14 118
rect -18 115 -14 116
rect -43 108 -42 110
rect -40 108 -39 110
rect -43 107 -39 108
rect -1 110 3 200
rect 74 202 78 203
rect 74 200 75 202
rect 77 200 78 202
rect 74 198 78 200
rect 74 196 75 198
rect 77 196 78 198
rect 74 195 78 196
rect 114 198 118 211
rect 347 213 351 214
rect 347 211 348 213
rect 350 211 351 213
rect 114 196 115 198
rect 117 196 118 198
rect 114 194 118 196
rect 303 202 307 203
rect 303 200 304 202
rect 306 200 307 202
rect 303 198 307 200
rect 303 196 304 198
rect 306 196 307 198
rect 303 194 307 196
rect 347 198 351 211
rect 347 196 348 198
rect 350 196 351 198
rect 347 194 351 196
rect 416 202 420 203
rect 416 200 417 202
rect 419 200 420 202
rect 416 198 420 200
rect 416 196 417 198
rect 419 196 420 198
rect 416 195 420 196
rect 460 202 464 204
rect 460 200 461 202
rect 463 200 464 202
rect 460 198 464 200
rect 460 196 461 198
rect 463 196 464 198
rect 460 194 464 196
rect 543 203 547 204
rect 543 201 544 203
rect 546 201 547 203
rect 543 197 547 201
rect 543 195 544 197
rect 546 195 547 197
rect 586 203 590 204
rect 586 201 587 203
rect 589 201 590 203
rect 586 198 590 201
rect 586 196 587 198
rect 589 196 590 198
rect 586 195 590 196
rect 669 203 673 204
rect 669 201 670 203
rect 672 201 673 203
rect 669 198 673 201
rect 669 196 670 198
rect 672 196 673 198
rect 669 195 673 196
rect 543 194 547 195
rect 157 193 161 194
rect 157 191 158 193
rect 160 191 161 193
rect 157 189 161 191
rect 157 187 158 189
rect 160 187 161 189
rect 157 186 161 187
rect 261 193 265 194
rect 261 191 262 193
rect 264 191 265 193
rect 261 189 265 191
rect 261 187 262 189
rect 264 187 265 189
rect 261 186 265 187
rect 502 193 506 194
rect 502 191 503 193
rect 505 191 506 193
rect 502 189 506 191
rect 502 187 503 189
rect 505 187 506 189
rect 502 186 506 187
rect 626 193 630 194
rect 626 191 627 193
rect 629 191 630 193
rect 626 189 630 191
rect 626 187 627 189
rect 629 187 630 189
rect 626 186 630 187
rect 66 180 71 182
rect 66 178 67 180
rect 69 178 71 180
rect 47 164 51 167
rect 47 162 48 164
rect 50 162 51 164
rect 47 126 51 162
rect 66 161 71 178
rect 106 181 111 182
rect 106 179 107 181
rect 109 179 111 181
rect 106 177 111 179
rect 106 175 108 177
rect 110 175 111 177
rect 295 181 300 182
rect 295 179 296 181
rect 298 179 300 181
rect 295 177 300 179
rect 295 175 297 177
rect 299 175 300 177
rect 106 174 111 175
rect 149 172 154 174
rect 149 170 151 172
rect 153 170 154 172
rect 66 159 67 161
rect 69 159 71 161
rect 66 158 71 159
rect 82 164 87 167
rect 82 162 84 164
rect 86 162 87 164
rect 47 124 48 126
rect 50 124 51 126
rect 47 122 51 124
rect 63 133 68 134
rect 63 131 65 133
rect 67 131 68 133
rect 63 119 68 131
rect 82 133 87 162
rect 126 164 130 167
rect 126 162 127 164
rect 129 162 130 164
rect 82 131 84 133
rect 86 131 87 133
rect 82 130 87 131
rect 114 132 118 133
rect 114 130 115 132
rect 117 130 118 132
rect 114 127 118 130
rect 114 125 115 127
rect 117 125 118 127
rect 114 124 118 125
rect 63 117 64 119
rect 66 117 68 119
rect 63 115 68 117
rect -1 108 0 110
rect 2 108 3 110
rect -1 107 3 108
rect -75 105 -71 106
rect -75 103 -74 105
rect -72 103 -71 105
rect -160 53 -159 55
rect -157 53 -156 55
rect -160 52 -156 53
rect -84 61 -80 62
rect -84 59 -83 61
rect -81 59 -80 61
rect -84 55 -80 59
rect -75 61 -71 103
rect -75 59 -74 61
rect -72 59 -71 61
rect -75 58 -71 59
rect -33 104 -28 106
rect -33 102 -32 104
rect -30 102 -28 104
rect -84 53 -83 55
rect -81 53 -80 55
rect -84 52 -80 53
rect -177 36 -176 38
rect -174 36 -173 38
rect -177 35 -173 36
rect -117 46 -112 47
rect -117 44 -115 46
rect -113 44 -112 46
rect -117 38 -112 44
rect -33 46 -28 102
rect -33 44 -32 46
rect -30 44 -28 46
rect -33 43 -28 44
rect 14 105 19 107
rect 14 103 16 105
rect 18 103 19 105
rect -117 36 -115 38
rect -113 36 -112 38
rect -117 34 -112 36
rect -11 35 -7 36
rect -11 33 -10 35
rect -8 33 -7 35
rect -108 30 -104 31
rect -140 29 -136 30
rect -140 27 -139 29
rect -137 27 -136 29
rect -140 24 -136 27
rect -192 21 -188 23
rect -140 22 -139 24
rect -137 22 -136 24
rect -192 19 -191 21
rect -189 19 -188 21
rect -202 -12 -198 -11
rect -202 -14 -201 -12
rect -199 -14 -198 -12
rect -202 -17 -198 -14
rect -202 -19 -201 -17
rect -199 -19 -198 -17
rect -202 -20 -198 -19
rect -192 -34 -188 19
rect -148 21 -144 22
rect -140 21 -136 22
rect -108 28 -107 30
rect -105 28 -104 30
rect -108 24 -104 28
rect -108 22 -107 24
rect -105 22 -104 24
rect -75 30 -71 31
rect -75 28 -74 30
rect -72 28 -71 30
rect -75 26 -71 28
rect -75 24 -74 26
rect -72 24 -71 26
rect -11 28 -7 33
rect -11 26 -10 28
rect -8 26 -7 28
rect -11 24 -7 26
rect 14 28 19 103
rect 114 102 118 104
rect 114 100 115 102
rect 117 100 118 102
rect 86 94 90 95
rect 86 92 87 94
rect 89 92 90 94
rect 53 61 57 62
rect 53 59 54 61
rect 56 59 57 61
rect 53 54 57 59
rect 53 52 54 54
rect 56 52 57 54
rect 53 51 57 52
rect 37 46 43 47
rect 37 44 39 46
rect 41 44 43 46
rect 37 37 43 44
rect 86 46 90 92
rect 114 61 118 100
rect 126 84 130 162
rect 149 150 154 170
rect 253 173 258 175
rect 295 174 300 175
rect 494 181 499 182
rect 494 179 495 181
rect 497 179 499 181
rect 494 177 499 179
rect 494 175 495 177
rect 497 175 499 177
rect 494 174 499 175
rect 578 181 583 182
rect 578 179 579 181
rect 581 179 583 181
rect 578 177 583 179
rect 578 175 579 177
rect 581 175 583 177
rect 578 174 583 175
rect 253 171 254 173
rect 256 171 258 173
rect 149 148 150 150
rect 152 148 154 150
rect 149 147 154 148
rect 233 164 237 167
rect 233 162 234 164
rect 236 162 237 164
rect 146 132 150 133
rect 146 130 147 132
rect 149 130 150 132
rect 146 126 150 130
rect 146 124 147 126
rect 149 124 150 126
rect 146 123 150 124
rect 179 130 183 131
rect 179 128 180 130
rect 182 128 183 130
rect 179 126 183 128
rect 233 130 237 162
rect 253 161 258 171
rect 315 173 319 174
rect 315 171 316 173
rect 318 171 319 173
rect 253 159 255 161
rect 257 159 258 161
rect 253 158 258 159
rect 271 164 275 167
rect 271 162 272 164
rect 274 162 275 164
rect 233 128 234 130
rect 236 128 237 130
rect 233 127 237 128
rect 243 128 247 130
rect 179 124 180 126
rect 182 124 183 126
rect 179 123 183 124
rect 243 126 244 128
rect 246 126 247 128
rect 243 121 247 126
rect 137 118 142 120
rect 243 119 244 121
rect 246 119 247 121
rect 243 118 247 119
rect 137 116 139 118
rect 141 116 142 118
rect 137 110 142 116
rect 137 108 139 110
rect 141 108 142 110
rect 137 107 142 108
rect 271 110 275 162
rect 271 108 272 110
rect 274 108 275 110
rect 271 107 275 108
rect 291 119 297 120
rect 291 117 292 119
rect 294 117 297 119
rect 291 110 297 117
rect 315 119 319 171
rect 339 173 344 174
rect 339 171 340 173
rect 342 171 344 173
rect 339 169 344 171
rect 339 167 340 169
rect 342 167 344 169
rect 408 173 413 174
rect 408 171 409 173
rect 411 171 413 173
rect 408 169 413 171
rect 408 167 409 169
rect 411 167 413 169
rect 339 166 344 167
rect 387 164 391 167
rect 408 166 413 167
rect 452 173 457 174
rect 452 171 453 173
rect 455 171 457 173
rect 387 162 388 164
rect 390 162 391 164
rect 332 132 336 133
rect 332 130 333 132
rect 335 130 336 132
rect 332 127 336 130
rect 332 125 333 127
rect 335 125 336 127
rect 332 124 336 125
rect 364 132 368 133
rect 364 130 365 132
rect 367 130 368 132
rect 364 126 368 130
rect 364 124 365 126
rect 367 124 368 126
rect 364 123 368 124
rect 387 126 391 162
rect 436 165 440 166
rect 436 163 437 165
rect 439 163 440 165
rect 387 124 388 126
rect 390 124 391 126
rect 387 122 391 124
rect 397 130 401 131
rect 397 128 398 130
rect 400 128 401 130
rect 397 126 401 128
rect 397 124 398 126
rect 400 124 401 126
rect 397 123 401 124
rect 315 117 316 119
rect 318 117 319 119
rect 315 116 319 117
rect 355 118 360 120
rect 355 116 357 118
rect 359 116 360 118
rect 291 108 293 110
rect 295 108 297 110
rect 291 107 297 108
rect 355 110 360 116
rect 355 108 357 110
rect 359 108 360 110
rect 355 107 360 108
rect 199 102 203 103
rect 170 101 174 102
rect 170 99 171 101
rect 173 99 174 101
rect 170 95 174 99
rect 170 93 171 95
rect 173 93 174 95
rect 170 92 174 93
rect 199 100 200 102
rect 202 100 203 102
rect 126 82 127 84
rect 129 82 130 84
rect 126 81 130 82
rect 143 84 147 89
rect 143 82 144 84
rect 146 82 147 84
rect 114 59 115 61
rect 117 59 118 61
rect 114 58 118 59
rect 134 61 138 62
rect 134 59 135 61
rect 137 59 138 61
rect 134 55 138 59
rect 134 53 135 55
rect 137 53 138 55
rect 134 52 138 53
rect 86 44 87 46
rect 89 44 90 46
rect 86 43 90 44
rect 101 46 106 47
rect 101 44 103 46
rect 105 44 106 46
rect 37 35 38 37
rect 40 35 43 37
rect 37 34 43 35
rect 101 38 106 44
rect 101 36 103 38
rect 105 36 106 38
rect 101 34 106 36
rect 110 30 114 31
rect 14 26 15 28
rect 17 26 19 28
rect 14 24 19 26
rect 78 29 82 30
rect 78 27 79 29
rect 81 27 82 29
rect 78 24 82 27
rect -75 23 -71 24
rect -108 21 -104 22
rect -48 22 -44 23
rect 78 22 79 24
rect 81 22 82 24
rect -148 19 -147 21
rect -145 19 -144 21
rect -170 -12 -166 -11
rect -170 -14 -169 -12
rect -167 -14 -166 -12
rect -170 -18 -166 -14
rect -148 -14 -144 19
rect -48 20 -47 22
rect -45 20 -44 22
rect -48 9 -44 20
rect 70 21 74 22
rect 78 21 82 22
rect 110 28 111 30
rect 113 28 114 30
rect 110 24 114 28
rect 110 22 111 24
rect 113 22 114 24
rect 143 30 147 82
rect 199 82 203 100
rect 307 102 311 103
rect 307 100 308 102
rect 310 100 311 102
rect 307 95 311 100
rect 307 93 308 95
rect 310 93 311 95
rect 307 92 311 93
rect 332 102 336 104
rect 420 102 424 103
rect 332 100 333 102
rect 335 100 336 102
rect 199 80 200 82
rect 202 80 203 82
rect 199 79 203 80
rect 321 82 326 83
rect 321 80 323 82
rect 325 80 326 82
rect 271 61 275 62
rect 271 59 272 61
rect 274 59 275 61
rect 271 54 275 59
rect 271 52 272 54
rect 274 52 275 54
rect 271 51 275 52
rect 255 46 261 47
rect 255 44 257 46
rect 259 44 261 46
rect 255 37 261 44
rect 143 28 144 30
rect 146 28 147 30
rect 143 26 147 28
rect 143 24 144 26
rect 146 24 147 26
rect 207 35 211 36
rect 207 33 208 35
rect 210 33 211 35
rect 255 35 256 37
rect 258 35 261 37
rect 255 34 261 35
rect 321 46 326 80
rect 332 61 336 100
rect 388 101 392 102
rect 388 99 389 101
rect 391 99 392 101
rect 388 95 392 99
rect 388 93 389 95
rect 391 93 392 95
rect 388 92 392 93
rect 420 100 421 102
rect 423 100 424 102
rect 420 84 424 100
rect 420 82 421 84
rect 423 82 424 84
rect 420 81 424 82
rect 332 59 333 61
rect 335 59 336 61
rect 332 58 336 59
rect 345 61 349 62
rect 345 59 346 61
rect 348 59 349 61
rect 321 44 323 46
rect 325 44 326 46
rect 321 38 326 44
rect 321 36 323 38
rect 325 36 326 38
rect 321 34 326 36
rect 345 38 349 59
rect 354 61 358 62
rect 354 59 355 61
rect 357 59 358 61
rect 354 55 358 59
rect 436 61 440 163
rect 452 151 457 171
rect 535 173 540 174
rect 535 171 536 173
rect 538 171 540 173
rect 452 149 453 151
rect 455 149 457 151
rect 452 147 457 149
rect 470 164 474 165
rect 470 162 471 164
rect 473 162 474 164
rect 461 128 465 130
rect 461 126 462 128
rect 464 126 465 128
rect 461 121 465 126
rect 461 119 462 121
rect 464 119 465 121
rect 461 118 465 119
rect 470 110 474 162
rect 518 164 523 166
rect 518 162 519 164
rect 521 162 523 164
rect 518 134 523 162
rect 535 161 540 171
rect 619 172 623 174
rect 619 170 620 172
rect 622 170 623 172
rect 619 169 623 170
rect 619 167 620 169
rect 622 167 623 169
rect 535 159 537 161
rect 539 159 540 161
rect 535 158 540 159
rect 561 164 566 167
rect 619 166 623 167
rect 662 172 666 174
rect 662 170 663 172
rect 665 170 666 172
rect 662 169 666 170
rect 662 167 663 169
rect 665 167 666 169
rect 662 166 666 167
rect 561 162 562 164
rect 564 162 566 164
rect 518 132 519 134
rect 521 132 523 134
rect 518 131 523 132
rect 533 134 537 135
rect 533 132 534 134
rect 536 132 537 134
rect 470 108 471 110
rect 473 108 474 110
rect 470 107 474 108
rect 509 119 515 120
rect 509 117 510 119
rect 512 117 515 119
rect 509 110 515 117
rect 533 119 537 132
rect 561 134 566 162
rect 601 164 606 165
rect 601 162 602 164
rect 604 162 606 164
rect 561 132 562 134
rect 564 132 566 134
rect 561 131 566 132
rect 585 134 589 135
rect 585 132 586 134
rect 588 132 589 134
rect 585 126 589 132
rect 585 124 586 126
rect 588 124 589 126
rect 585 123 589 124
rect 533 117 534 119
rect 536 117 537 119
rect 533 116 537 117
rect 601 119 606 162
rect 601 117 602 119
rect 604 117 606 119
rect 601 116 606 117
rect 509 108 511 110
rect 513 108 515 110
rect 509 107 515 108
rect 552 106 558 111
rect 552 104 554 106
rect 556 104 558 106
rect 525 102 529 103
rect 525 100 526 102
rect 528 100 529 102
rect 525 95 529 100
rect 525 93 526 95
rect 528 93 529 95
rect 525 92 529 93
rect 535 84 539 85
rect 535 82 536 84
rect 538 82 539 84
rect 436 59 437 61
rect 439 59 440 61
rect 436 58 440 59
rect 491 61 495 62
rect 491 59 492 61
rect 494 59 495 61
rect 354 53 355 55
rect 357 53 358 55
rect 354 52 358 53
rect 491 54 495 59
rect 491 52 492 54
rect 494 52 495 54
rect 491 51 495 52
rect 345 36 346 38
rect 348 36 349 38
rect 475 46 481 47
rect 475 44 477 46
rect 479 44 481 46
rect 475 37 481 44
rect 345 35 349 36
rect 427 35 431 36
rect 207 28 211 33
rect 427 33 428 35
rect 430 33 431 35
rect 475 35 476 37
rect 478 35 481 37
rect 535 38 539 82
rect 552 46 558 104
rect 552 44 553 46
rect 555 44 558 46
rect 552 43 558 44
rect 535 36 536 38
rect 538 36 539 38
rect 535 35 539 36
rect 475 34 481 35
rect 330 30 334 31
rect 207 26 208 28
rect 210 26 211 28
rect 207 24 211 26
rect 298 29 302 30
rect 298 27 299 29
rect 301 27 302 29
rect 298 24 302 27
rect 143 23 147 24
rect 110 21 114 22
rect 169 22 173 23
rect 298 22 299 24
rect 301 22 302 24
rect 70 19 71 21
rect 73 19 74 21
rect -48 7 -47 9
rect -45 7 -44 9
rect -48 6 -44 7
rect 41 9 46 10
rect 41 7 43 9
rect 45 7 46 9
rect 18 -12 22 -11
rect -148 -16 -147 -14
rect -145 -16 -144 -14
rect -148 -17 -144 -16
rect -137 -14 -133 -13
rect 18 -14 19 -12
rect 21 -14 22 -12
rect -137 -16 -136 -14
rect -134 -16 -133 -14
rect -170 -20 -169 -18
rect -167 -20 -166 -18
rect -170 -21 -166 -20
rect -137 -18 -133 -16
rect -137 -20 -136 -18
rect -134 -20 -133 -18
rect -137 -21 -133 -20
rect -73 -16 -69 -14
rect -73 -18 -72 -16
rect -70 -18 -69 -16
rect -73 -23 -69 -18
rect 18 -17 22 -14
rect 18 -19 19 -17
rect 21 -19 22 -17
rect 18 -20 22 -19
rect -192 -36 -191 -34
rect -189 -36 -188 -34
rect -192 -37 -188 -36
rect -179 -26 -174 -24
rect -73 -25 -72 -23
rect -70 -25 -69 -23
rect -73 -26 -69 -25
rect -25 -25 -19 -24
rect -179 -28 -177 -26
rect -175 -28 -174 -26
rect -179 -34 -174 -28
rect -179 -36 -177 -34
rect -175 -36 -174 -34
rect -179 -37 -174 -36
rect -25 -27 -24 -25
rect -22 -27 -19 -25
rect -25 -34 -19 -27
rect -25 -36 -23 -34
rect -21 -36 -19 -34
rect -25 -37 -19 -36
rect 41 -26 46 7
rect 50 -12 54 -11
rect 50 -14 51 -12
rect 53 -14 54 -12
rect 50 -18 54 -14
rect 70 -14 74 19
rect 169 20 170 22
rect 172 20 173 22
rect 169 9 173 20
rect 290 21 294 22
rect 298 21 302 22
rect 330 28 331 30
rect 333 28 334 30
rect 330 24 334 28
rect 330 22 331 24
rect 333 22 334 24
rect 363 30 367 31
rect 363 28 364 30
rect 366 28 367 30
rect 363 26 367 28
rect 363 24 364 26
rect 366 24 367 26
rect 427 28 431 33
rect 427 26 428 28
rect 430 26 431 28
rect 427 24 431 26
rect 511 25 515 27
rect 363 23 367 24
rect 511 23 512 25
rect 514 23 515 25
rect 330 21 334 22
rect 390 22 394 23
rect 290 19 291 21
rect 293 19 294 21
rect 169 7 170 9
rect 172 7 173 9
rect 169 6 173 7
rect 258 9 263 10
rect 258 7 259 9
rect 261 7 263 9
rect 235 -12 239 -11
rect 70 -16 71 -14
rect 73 -16 74 -14
rect 70 -17 74 -16
rect 83 -14 87 -13
rect 235 -14 236 -12
rect 238 -14 239 -12
rect 83 -16 84 -14
rect 86 -16 87 -14
rect 50 -20 51 -18
rect 53 -20 54 -18
rect 50 -21 54 -20
rect 83 -18 87 -16
rect 83 -20 84 -18
rect 86 -20 87 -18
rect 83 -21 87 -20
rect 147 -16 151 -14
rect 147 -18 148 -16
rect 150 -18 151 -16
rect 147 -23 151 -18
rect 235 -17 239 -14
rect 235 -19 236 -17
rect 238 -19 239 -17
rect 235 -20 239 -19
rect 147 -25 148 -23
rect 150 -25 151 -23
rect 147 -26 151 -25
rect 195 -25 201 -24
rect 41 -28 43 -26
rect 45 -28 46 -26
rect 41 -34 46 -28
rect 41 -36 43 -34
rect 45 -36 46 -34
rect 41 -37 46 -36
rect 195 -27 196 -25
rect 198 -27 201 -25
rect 195 -34 201 -27
rect 195 -36 197 -34
rect 199 -36 201 -34
rect 195 -37 201 -36
rect 258 -26 263 7
rect 267 -12 271 -11
rect 267 -14 268 -12
rect 270 -14 271 -12
rect 267 -18 271 -14
rect 267 -20 268 -18
rect 270 -20 271 -18
rect 267 -21 271 -20
rect 290 -18 294 19
rect 390 20 391 22
rect 393 20 394 22
rect 390 9 394 20
rect 390 7 391 9
rect 393 7 394 9
rect 390 6 394 7
rect 470 9 475 10
rect 470 7 471 9
rect 473 7 475 9
rect 290 -20 291 -18
rect 293 -20 294 -18
rect 290 -21 294 -20
rect 300 -14 304 -13
rect 300 -16 301 -14
rect 303 -16 304 -14
rect 300 -18 304 -16
rect 300 -20 301 -18
rect 303 -20 304 -18
rect 300 -21 304 -20
rect 364 -16 368 -14
rect 364 -18 365 -16
rect 367 -18 368 -16
rect 364 -23 368 -18
rect 364 -25 365 -23
rect 367 -25 368 -23
rect 364 -26 368 -25
rect 412 -25 418 -24
rect 258 -28 260 -26
rect 262 -28 263 -26
rect 258 -34 263 -28
rect 258 -36 260 -34
rect 262 -36 263 -34
rect 258 -37 263 -36
rect 412 -27 413 -25
rect 415 -27 418 -25
rect 412 -34 418 -27
rect 412 -36 414 -34
rect 416 -36 418 -34
rect 412 -37 418 -36
rect 470 -34 475 7
rect 487 9 491 10
rect 487 7 488 9
rect 490 7 491 9
rect 487 -17 491 7
rect 511 9 515 23
rect 511 7 512 9
rect 514 7 515 9
rect 511 6 515 7
rect 487 -19 488 -17
rect 490 -19 491 -17
rect 487 -20 491 -19
rect 470 -36 472 -34
rect 474 -36 475 -34
rect 470 -37 475 -36
rect 10 -39 14 -37
rect 10 -41 11 -39
rect 13 -41 14 -39
rect 227 -38 231 -37
rect 227 -40 228 -38
rect 230 -40 231 -38
rect -9 -42 -5 -41
rect -146 -43 -142 -42
rect -146 -45 -145 -43
rect -143 -45 -142 -43
rect -146 -49 -142 -45
rect -146 -51 -145 -49
rect -143 -51 -142 -49
rect -146 -52 -142 -51
rect -9 -44 -8 -42
rect -6 -44 -5 -42
rect -9 -49 -5 -44
rect -9 -51 -8 -49
rect -6 -51 -5 -49
rect -9 -52 -5 -51
rect 10 -49 14 -41
rect 211 -42 215 -41
rect 10 -51 11 -49
rect 13 -51 14 -49
rect 10 -52 14 -51
rect 74 -43 78 -42
rect 74 -45 75 -43
rect 77 -45 78 -43
rect 74 -49 78 -45
rect 74 -51 75 -49
rect 77 -51 78 -49
rect 74 -52 78 -51
rect 211 -44 212 -42
rect 214 -44 215 -42
rect 211 -49 215 -44
rect 211 -51 212 -49
rect 214 -51 215 -49
rect 211 -52 215 -51
rect 227 -49 231 -40
rect 454 -39 458 -38
rect 454 -41 455 -39
rect 457 -41 458 -39
rect 428 -42 432 -41
rect 227 -51 228 -49
rect 230 -51 231 -49
rect 227 -52 231 -51
rect 291 -43 295 -42
rect 291 -45 292 -43
rect 294 -45 295 -43
rect 291 -49 295 -45
rect 291 -51 292 -49
rect 294 -51 295 -49
rect 291 -52 295 -51
rect 428 -44 429 -42
rect 431 -44 432 -42
rect 428 -49 432 -44
rect 428 -51 429 -49
rect 431 -51 432 -49
rect 428 -52 432 -51
rect 454 -49 458 -41
rect 454 -51 455 -49
rect 457 -51 458 -49
rect 454 -52 458 -51
<< alu3 >>
rect -160 213 351 214
rect -160 211 -159 213
rect -157 211 -42 213
rect -40 211 115 213
rect 117 211 348 213
rect 350 211 351 213
rect -160 210 351 211
rect 460 203 673 204
rect -1 202 420 203
rect -1 200 0 202
rect 2 200 75 202
rect 77 200 304 202
rect 306 200 417 202
rect 419 200 420 202
rect -1 199 420 200
rect 460 202 544 203
rect 460 200 461 202
rect 463 201 544 202
rect 546 201 587 203
rect 589 201 670 203
rect 672 201 673 203
rect 463 200 673 201
rect 460 199 673 200
rect 157 189 630 190
rect 157 187 158 189
rect 160 187 262 189
rect 264 187 503 189
rect 505 187 627 189
rect 629 187 630 189
rect 157 186 630 187
rect 106 177 583 178
rect 106 175 108 177
rect 110 175 297 177
rect 299 175 495 177
rect 497 175 579 177
rect 581 175 583 177
rect 106 174 583 175
rect 339 169 666 170
rect 339 167 340 169
rect 342 167 409 169
rect 411 167 620 169
rect 622 167 663 169
rect 665 167 666 169
rect 339 166 666 167
rect -60 161 540 162
rect -60 159 -59 161
rect -57 159 67 161
rect 69 159 255 161
rect 257 159 537 161
rect 539 159 540 161
rect -60 158 540 159
rect -177 151 457 152
rect -177 150 453 151
rect -177 148 -176 150
rect -174 148 -17 150
rect -15 148 150 150
rect 152 149 453 150
rect 455 149 457 151
rect 152 148 457 149
rect -177 147 457 148
rect 518 134 537 135
rect 63 133 87 134
rect 63 131 65 133
rect 67 131 84 133
rect 86 131 87 133
rect 63 130 87 131
rect 114 132 151 133
rect 114 130 115 132
rect 117 130 147 132
rect 149 130 151 132
rect 332 132 369 133
rect 114 129 151 130
rect 179 130 247 131
rect 179 128 180 130
rect 182 128 234 130
rect 236 128 247 130
rect 332 130 333 132
rect 335 130 365 132
rect 367 130 369 132
rect 518 132 519 134
rect 521 132 534 134
rect 536 132 537 134
rect 518 131 537 132
rect 561 134 589 135
rect 561 132 562 134
rect 564 132 586 134
rect 588 132 589 134
rect 561 131 589 132
rect 332 129 369 130
rect 397 130 465 131
rect 179 127 244 128
rect 243 126 244 127
rect 246 126 247 128
rect 397 128 398 130
rect 400 128 465 130
rect 397 127 462 128
rect 243 125 247 126
rect 461 126 462 127
rect 464 126 465 128
rect 461 125 465 126
rect 137 110 297 111
rect 137 108 139 110
rect 141 108 272 110
rect 274 108 293 110
rect 295 108 297 110
rect 137 107 297 108
rect 355 110 515 111
rect 355 108 357 110
rect 359 108 471 110
rect 473 108 511 110
rect 513 108 515 110
rect 355 107 515 108
rect 170 95 311 96
rect 170 93 171 95
rect 173 93 308 95
rect 310 93 311 95
rect 170 92 311 93
rect 388 95 529 96
rect 388 93 389 95
rect 391 93 526 95
rect 528 93 529 95
rect 388 92 529 93
rect 126 84 147 85
rect 126 82 127 84
rect 129 82 144 84
rect 146 82 147 84
rect 420 84 539 85
rect 126 81 147 82
rect 199 82 326 83
rect 199 80 200 82
rect 202 80 323 82
rect 325 80 326 82
rect 420 82 421 84
rect 423 82 536 84
rect 538 82 539 84
rect 420 81 539 82
rect 199 79 326 80
rect -84 61 57 62
rect -84 59 -83 61
rect -81 59 -74 61
rect -72 59 54 61
rect 56 59 57 61
rect -84 58 57 59
rect 114 61 275 62
rect 114 59 115 61
rect 117 59 135 61
rect 137 59 272 61
rect 274 59 275 61
rect 114 58 275 59
rect 332 61 349 62
rect 332 59 333 61
rect 335 59 346 61
rect 348 59 349 61
rect 332 58 349 59
rect 354 61 495 62
rect 354 59 355 61
rect 357 59 437 61
rect 439 59 492 61
rect 494 59 495 61
rect 354 58 495 59
rect -117 46 43 47
rect -117 44 -115 46
rect -113 44 -32 46
rect -30 44 39 46
rect 41 44 43 46
rect -117 43 43 44
rect 86 46 261 47
rect 86 44 87 46
rect 89 44 103 46
rect 105 44 257 46
rect 259 44 261 46
rect 86 43 261 44
rect 321 46 481 47
rect 321 44 323 46
rect 325 44 477 46
rect 479 44 481 46
rect 321 43 481 44
rect -11 28 19 29
rect -11 27 -10 28
rect -75 26 -10 27
rect -8 26 15 28
rect 17 26 19 28
rect 207 28 211 29
rect 207 27 208 28
rect -140 24 -103 25
rect -140 22 -139 24
rect -137 22 -107 24
rect -105 22 -103 24
rect -75 24 -74 26
rect -72 24 19 26
rect 143 26 208 27
rect 210 26 211 28
rect 427 28 431 29
rect 427 27 428 28
rect 78 24 115 25
rect -75 23 -7 24
rect -140 21 -103 22
rect 78 22 79 24
rect 81 22 111 24
rect 113 22 115 24
rect 143 24 144 26
rect 146 24 211 26
rect 363 26 428 27
rect 430 26 431 28
rect 143 23 211 24
rect 298 24 335 25
rect 78 21 115 22
rect 298 22 299 24
rect 301 22 331 24
rect 333 22 335 24
rect 363 24 364 26
rect 366 24 431 26
rect 363 23 431 24
rect 298 21 335 22
rect -48 9 46 10
rect -48 7 -47 9
rect -45 7 43 9
rect 45 7 46 9
rect -48 6 46 7
rect 169 9 263 10
rect 169 7 170 9
rect 172 7 259 9
rect 261 7 263 9
rect 169 6 263 7
rect 390 9 475 10
rect 390 7 391 9
rect 393 7 471 9
rect 473 7 475 9
rect 390 6 475 7
rect 487 9 515 10
rect 487 7 488 9
rect 490 7 512 9
rect 514 7 515 9
rect 487 6 515 7
rect -202 -12 -165 -11
rect -202 -14 -201 -12
rect -199 -14 -169 -12
rect -167 -14 -165 -12
rect 18 -12 55 -11
rect -202 -15 -165 -14
rect -148 -14 -69 -13
rect -148 -16 -147 -14
rect -145 -16 -136 -14
rect -134 -16 -69 -14
rect 18 -14 19 -12
rect 21 -14 51 -12
rect 53 -14 55 -12
rect 235 -12 272 -11
rect 18 -15 55 -14
rect 70 -14 151 -13
rect -148 -17 -72 -16
rect -73 -18 -72 -17
rect -70 -18 -69 -16
rect 70 -16 71 -14
rect 73 -16 84 -14
rect 86 -16 151 -14
rect 235 -14 236 -12
rect 238 -14 268 -12
rect 270 -14 272 -12
rect 235 -15 272 -14
rect 300 -14 368 -13
rect 70 -17 148 -16
rect -73 -19 -69 -18
rect 147 -18 148 -17
rect 150 -18 151 -16
rect 300 -16 301 -14
rect 303 -16 368 -14
rect 300 -17 365 -16
rect 147 -19 151 -18
rect 364 -18 365 -17
rect 367 -18 368 -16
rect 364 -19 368 -18
rect -192 -34 -19 -33
rect -192 -36 -191 -34
rect -189 -36 -177 -34
rect -175 -36 -23 -34
rect -21 -36 -19 -34
rect -192 -37 -19 -36
rect 41 -34 201 -33
rect 41 -36 43 -34
rect 45 -36 197 -34
rect 199 -36 201 -34
rect 41 -37 201 -36
rect 258 -34 418 -33
rect 258 -36 260 -34
rect 262 -36 414 -34
rect 416 -36 418 -34
rect 258 -37 418 -36
rect -146 -49 14 -48
rect -146 -51 -145 -49
rect -143 -51 -8 -49
rect -6 -51 11 -49
rect 13 -51 14 -49
rect -146 -52 14 -51
rect 74 -49 231 -48
rect 74 -51 75 -49
rect 77 -51 212 -49
rect 214 -51 228 -49
rect 230 -51 231 -49
rect 74 -52 231 -51
rect 291 -49 458 -48
rect 291 -51 292 -49
rect 294 -51 429 -49
rect 431 -51 455 -49
rect 457 -51 458 -49
rect 291 -52 458 -51
<< ptie >>
rect 43 155 49 157
rect 43 153 45 155
rect 47 153 49 155
rect 43 151 49 153
rect 83 155 89 157
rect 83 153 85 155
rect 87 153 89 155
rect 83 151 89 153
rect 126 155 132 157
rect 126 153 128 155
rect 130 153 132 155
rect 126 151 132 153
rect 230 155 236 157
rect 230 153 232 155
rect 234 153 236 155
rect 230 151 236 153
rect 272 155 278 157
rect 272 153 274 155
rect 276 153 278 155
rect 272 151 278 153
rect 316 155 322 157
rect 316 153 318 155
rect 320 153 322 155
rect 316 151 322 153
rect 385 155 391 157
rect 385 153 387 155
rect 389 153 391 155
rect 385 151 391 153
rect 429 155 435 157
rect 429 153 431 155
rect 433 153 435 155
rect 429 151 435 153
rect 471 155 477 157
rect 471 153 473 155
rect 475 153 477 155
rect 471 151 477 153
rect 512 155 518 157
rect 512 153 514 155
rect 516 153 518 155
rect 512 151 518 153
rect 555 155 561 157
rect 555 153 557 155
rect 559 153 561 155
rect 555 151 561 153
rect 595 155 601 157
rect 595 153 597 155
rect 599 153 601 155
rect 595 151 601 153
rect 638 155 644 157
rect 638 153 640 155
rect 642 153 644 155
rect 638 151 644 153
rect -74 144 -68 146
rect -74 142 -72 144
rect -70 142 -68 144
rect -74 140 -68 142
rect -32 144 -26 146
rect -32 142 -30 144
rect -28 142 -26 144
rect -32 140 -26 142
rect 107 144 125 146
rect 107 142 109 144
rect 111 142 121 144
rect 123 142 125 144
rect 107 140 125 142
rect 312 144 318 146
rect 312 142 314 144
rect 316 142 318 144
rect 312 140 318 142
rect 325 144 343 146
rect 325 142 327 144
rect 329 142 339 144
rect 341 142 343 144
rect 325 140 343 142
rect 530 144 536 146
rect 530 142 532 144
rect 534 142 536 144
rect 530 140 536 142
rect -191 12 -185 14
rect -191 10 -189 12
rect -187 10 -185 12
rect -191 8 -185 10
rect -147 12 -129 14
rect -147 10 -145 12
rect -143 10 -133 12
rect -131 10 -129 12
rect -147 8 -129 10
rect 58 12 64 14
rect 58 10 60 12
rect 62 10 64 12
rect 58 8 64 10
rect 71 12 89 14
rect 71 10 73 12
rect 75 10 85 12
rect 87 10 89 12
rect 71 8 89 10
rect 276 12 282 14
rect 276 10 278 12
rect 280 10 282 12
rect 276 8 282 10
rect 291 12 309 14
rect 291 10 293 12
rect 295 10 305 12
rect 307 10 309 12
rect 291 8 309 10
rect 496 12 502 14
rect 496 10 498 12
rect 500 10 502 12
rect 496 8 502 10
rect -209 0 -191 2
rect -209 -2 -207 0
rect -205 -2 -195 0
rect -193 -2 -191 0
rect -209 -4 -191 -2
rect -4 0 2 2
rect -4 -2 -2 0
rect 0 -2 2 0
rect -4 -4 2 -2
rect 11 0 29 2
rect 11 -2 13 0
rect 15 -2 25 0
rect 27 -2 29 0
rect 11 -4 29 -2
rect 216 0 222 2
rect 216 -2 218 0
rect 220 -2 222 0
rect 216 -4 222 -2
rect 228 0 246 2
rect 228 -2 230 0
rect 232 -2 242 0
rect 244 -2 246 0
rect 228 -4 246 -2
rect 433 0 439 2
rect 433 -2 435 0
rect 437 -2 439 0
rect 433 -4 439 -2
<< ntie >>
rect 43 215 49 217
rect 43 213 45 215
rect 47 213 49 215
rect 43 211 49 213
rect 83 215 89 217
rect 83 213 85 215
rect 87 213 89 215
rect 83 211 89 213
rect 126 215 132 217
rect 126 213 128 215
rect 130 213 132 215
rect 126 211 132 213
rect 230 215 236 217
rect 230 213 232 215
rect 234 213 236 215
rect 230 211 236 213
rect 272 215 278 217
rect 272 213 274 215
rect 276 213 278 215
rect 272 211 278 213
rect 316 215 322 217
rect 316 213 318 215
rect 320 213 322 215
rect 316 211 322 213
rect 385 215 391 217
rect 385 213 387 215
rect 389 213 391 215
rect 385 211 391 213
rect 429 215 435 217
rect 429 213 431 215
rect 433 213 435 215
rect 429 211 435 213
rect 471 215 477 217
rect 471 213 473 215
rect 475 213 477 215
rect 471 211 477 213
rect 512 215 518 217
rect 512 213 514 215
rect 516 213 518 215
rect 512 211 518 213
rect 555 215 561 217
rect 555 213 557 215
rect 559 213 561 215
rect 555 211 561 213
rect 595 215 601 217
rect 595 213 597 215
rect 599 213 601 215
rect 595 211 601 213
rect 638 215 644 217
rect 638 213 640 215
rect 642 213 644 215
rect 638 211 644 213
rect -74 84 -68 86
rect -74 82 -72 84
rect -70 82 -68 84
rect -74 80 -68 82
rect -32 84 -26 86
rect -32 82 -30 84
rect -28 82 -26 84
rect -32 80 -26 82
rect 107 84 125 86
rect 107 82 109 84
rect 111 82 121 84
rect 123 82 125 84
rect 107 80 125 82
rect 312 84 318 86
rect 312 82 314 84
rect 316 82 318 84
rect 312 80 318 82
rect 325 84 343 86
rect 325 82 327 84
rect 329 82 339 84
rect 341 82 343 84
rect 325 80 343 82
rect 530 84 536 86
rect 530 82 532 84
rect 534 82 536 84
rect 530 80 536 82
rect -191 72 -185 74
rect -191 70 -189 72
rect -187 70 -185 72
rect -191 68 -185 70
rect -147 72 -129 74
rect -147 70 -145 72
rect -143 70 -133 72
rect -131 70 -129 72
rect 58 72 64 74
rect -147 68 -129 70
rect 58 70 60 72
rect 62 70 64 72
rect 58 68 64 70
rect 71 72 89 74
rect 71 70 73 72
rect 75 70 85 72
rect 87 70 89 72
rect 276 72 282 74
rect 71 68 89 70
rect 276 70 278 72
rect 280 70 282 72
rect 276 68 282 70
rect 291 72 309 74
rect 291 70 293 72
rect 295 70 305 72
rect 307 70 309 72
rect 496 72 502 74
rect 291 68 309 70
rect 496 70 498 72
rect 500 70 502 72
rect 496 68 502 70
rect -209 -60 -191 -58
rect -209 -62 -207 -60
rect -205 -62 -195 -60
rect -193 -62 -191 -60
rect -209 -64 -191 -62
rect -4 -60 2 -58
rect -4 -62 -2 -60
rect 0 -62 2 -60
rect -4 -64 2 -62
rect 11 -60 29 -58
rect 11 -62 13 -60
rect 15 -62 25 -60
rect 27 -62 29 -60
rect 11 -64 29 -62
rect 216 -60 222 -58
rect 216 -62 218 -60
rect 220 -62 222 -60
rect 216 -64 222 -62
rect 228 -60 246 -58
rect 228 -62 230 -60
rect 232 -62 242 -60
rect 244 -62 246 -60
rect 228 -64 246 -62
rect 433 -60 439 -58
rect 433 -62 435 -60
rect 437 -62 439 -60
rect 433 -64 439 -62
<< nmos >>
rect 49 163 51 172
rect 62 161 64 172
rect 69 161 71 172
rect 89 163 91 172
rect 102 161 104 172
rect 109 161 111 172
rect 132 163 134 172
rect 145 161 147 172
rect 152 161 154 172
rect 236 163 238 172
rect 249 161 251 172
rect 256 161 258 172
rect 278 163 280 172
rect 291 161 293 172
rect 298 161 300 172
rect 322 163 324 172
rect 335 161 337 172
rect 342 161 344 172
rect 391 163 393 172
rect 404 161 406 172
rect 411 161 413 172
rect 435 163 437 172
rect 448 161 450 172
rect 455 161 457 172
rect 477 163 479 172
rect 490 161 492 172
rect 497 161 499 172
rect 518 163 520 172
rect 531 161 533 172
rect 538 161 540 172
rect 561 163 563 172
rect 574 161 576 172
rect 581 161 583 172
rect 601 163 603 172
rect 614 161 616 172
rect 621 161 623 172
rect 644 163 646 172
rect 657 161 659 172
rect 664 161 666 172
rect -68 125 -66 134
rect -55 125 -53 136
rect -48 125 -46 136
rect -26 125 -24 134
rect -13 125 -11 136
rect -6 125 -4 136
rect 22 129 24 143
rect 33 123 35 143
rect 40 123 42 143
rect 60 123 62 137
rect 70 123 72 137
rect 80 130 82 140
rect 90 130 92 143
rect 113 123 115 132
rect 137 125 139 137
rect 149 123 151 135
rect 156 123 158 135
rect 166 123 168 135
rect 176 123 178 135
rect 203 129 205 142
rect 210 129 212 142
rect 220 129 222 142
rect 230 124 232 137
rect 242 129 244 140
rect 265 129 267 142
rect 272 129 274 142
rect 282 129 284 142
rect 292 124 294 137
rect 303 123 305 134
rect 331 123 333 132
rect 355 125 357 137
rect 367 123 369 135
rect 374 123 376 135
rect 384 123 386 135
rect 394 123 396 135
rect 421 129 423 142
rect 428 129 430 142
rect 438 129 440 142
rect 448 124 450 137
rect 460 129 462 140
rect 483 129 485 142
rect 490 129 492 142
rect 500 129 502 142
rect 510 124 512 137
rect 521 123 523 134
rect 560 129 562 143
rect 571 123 573 143
rect 578 123 580 143
rect 598 123 600 137
rect 608 123 610 137
rect 618 130 620 140
rect 628 130 630 143
rect -185 20 -183 29
rect -172 18 -170 29
rect -165 18 -163 29
rect -141 22 -139 31
rect -117 17 -115 29
rect -105 19 -103 31
rect -98 19 -96 31
rect -88 19 -86 31
rect -78 19 -76 31
rect -51 12 -49 25
rect -44 12 -42 25
rect -34 12 -32 25
rect -24 17 -22 30
rect -12 14 -10 25
rect 11 12 13 25
rect 18 12 20 25
rect 28 12 30 25
rect 38 17 40 30
rect 49 20 51 31
rect 77 22 79 31
rect 101 17 103 29
rect 113 19 115 31
rect 120 19 122 31
rect 130 19 132 31
rect 140 19 142 31
rect 167 12 169 25
rect 174 12 176 25
rect 184 12 186 25
rect 194 17 196 30
rect 206 14 208 25
rect 229 12 231 25
rect 236 12 238 25
rect 246 12 248 25
rect 256 17 258 30
rect 267 20 269 31
rect 297 22 299 31
rect 321 17 323 29
rect 333 19 335 31
rect 340 19 342 31
rect 350 19 352 31
rect 360 19 362 31
rect 387 12 389 25
rect 394 12 396 25
rect 404 12 406 25
rect 414 17 416 30
rect 426 14 428 25
rect 449 12 451 25
rect 456 12 458 25
rect 466 12 468 25
rect 476 17 478 30
rect 487 20 489 31
rect 519 11 521 25
rect 530 11 532 31
rect 537 11 539 31
rect 557 17 559 31
rect 567 17 569 31
rect 577 14 579 24
rect 587 11 589 24
rect -203 -21 -201 -12
rect -179 -19 -177 -7
rect -167 -21 -165 -9
rect -160 -21 -158 -9
rect -150 -21 -148 -9
rect -140 -21 -138 -9
rect -113 -15 -111 -2
rect -106 -15 -104 -2
rect -96 -15 -94 -2
rect -86 -20 -84 -7
rect -74 -15 -72 -4
rect -51 -15 -49 -2
rect -44 -15 -42 -2
rect -34 -15 -32 -2
rect -24 -20 -22 -7
rect -13 -21 -11 -10
rect 17 -21 19 -12
rect 41 -19 43 -7
rect 53 -21 55 -9
rect 60 -21 62 -9
rect 70 -21 72 -9
rect 80 -21 82 -9
rect 107 -15 109 -2
rect 114 -15 116 -2
rect 124 -15 126 -2
rect 134 -20 136 -7
rect 146 -15 148 -4
rect 169 -15 171 -2
rect 176 -15 178 -2
rect 186 -15 188 -2
rect 196 -20 198 -7
rect 207 -21 209 -10
rect 234 -21 236 -12
rect 258 -19 260 -7
rect 270 -21 272 -9
rect 277 -21 279 -9
rect 287 -21 289 -9
rect 297 -21 299 -9
rect 324 -15 326 -2
rect 331 -15 333 -2
rect 341 -15 343 -2
rect 351 -20 353 -7
rect 363 -15 365 -4
rect 386 -15 388 -2
rect 393 -15 395 -2
rect 403 -15 405 -2
rect 413 -20 415 -7
rect 424 -21 426 -10
rect 462 -15 464 -1
rect 473 -21 475 -1
rect 480 -21 482 -1
rect 500 -21 502 -7
rect 510 -21 512 -7
rect 520 -14 522 -4
rect 530 -14 532 -1
<< pmos >>
rect 49 187 51 205
rect 59 194 61 207
rect 69 194 71 207
rect 89 187 91 205
rect 99 194 101 207
rect 109 194 111 207
rect 132 187 134 205
rect 142 194 144 207
rect 152 194 154 207
rect 236 187 238 205
rect 246 194 248 207
rect 256 194 258 207
rect 278 187 280 205
rect 288 194 290 207
rect 298 194 300 207
rect 322 187 324 205
rect 332 194 334 207
rect 342 194 344 207
rect 391 187 393 205
rect 401 194 403 207
rect 411 194 413 207
rect 435 187 437 205
rect 445 194 447 207
rect 455 194 457 207
rect 477 187 479 205
rect 487 194 489 207
rect 497 194 499 207
rect 518 187 520 205
rect 528 194 530 207
rect 538 194 540 207
rect 561 187 563 205
rect 571 194 573 207
rect 581 194 583 207
rect 601 187 603 205
rect 611 194 613 207
rect 621 194 623 207
rect 644 187 646 205
rect 654 194 656 207
rect 664 194 666 207
rect -68 92 -66 110
rect -58 90 -56 103
rect -48 90 -46 103
rect -26 92 -24 110
rect -16 90 -14 103
rect -6 90 -4 103
rect 22 83 24 111
rect 32 83 34 111
rect 42 83 44 111
rect 60 86 62 111
rect 67 86 69 111
rect 77 95 79 108
rect 90 83 92 108
rect 113 93 115 111
rect 140 84 142 111
rect 150 84 152 111
rect 157 84 159 111
rect 167 84 169 111
rect 177 84 179 111
rect 202 83 204 111
rect 212 83 214 111
rect 222 83 224 111
rect 232 83 234 97
rect 242 83 244 97
rect 262 83 264 111
rect 272 83 274 111
rect 282 83 284 111
rect 293 90 295 104
rect 303 90 305 104
rect 331 93 333 111
rect 358 84 360 111
rect 368 84 370 111
rect 375 84 377 111
rect 385 84 387 111
rect 395 84 397 111
rect 420 83 422 111
rect 430 83 432 111
rect 440 83 442 111
rect 450 83 452 97
rect 460 83 462 97
rect 480 83 482 111
rect 490 83 492 111
rect 500 83 502 111
rect 511 90 513 104
rect 521 90 523 104
rect 560 83 562 111
rect 570 83 572 111
rect 580 83 582 111
rect 598 86 600 111
rect 605 86 607 111
rect 615 95 617 108
rect 628 83 630 108
rect -185 44 -183 62
rect -175 51 -173 64
rect -165 51 -163 64
rect -141 43 -139 61
rect -114 43 -112 70
rect -104 43 -102 70
rect -97 43 -95 70
rect -87 43 -85 70
rect -77 43 -75 70
rect -52 43 -50 71
rect -42 43 -40 71
rect -32 43 -30 71
rect -22 57 -20 71
rect -12 57 -10 71
rect 8 43 10 71
rect 18 43 20 71
rect 28 43 30 71
rect 39 50 41 64
rect 49 50 51 64
rect 77 43 79 61
rect 104 43 106 70
rect 114 43 116 70
rect 121 43 123 70
rect 131 43 133 70
rect 141 43 143 70
rect 166 43 168 71
rect 176 43 178 71
rect 186 43 188 71
rect 196 57 198 71
rect 206 57 208 71
rect 226 43 228 71
rect 236 43 238 71
rect 246 43 248 71
rect 257 50 259 64
rect 267 50 269 64
rect 297 43 299 61
rect 324 43 326 70
rect 334 43 336 70
rect 341 43 343 70
rect 351 43 353 70
rect 361 43 363 70
rect 386 43 388 71
rect 396 43 398 71
rect 406 43 408 71
rect 416 57 418 71
rect 426 57 428 71
rect 446 43 448 71
rect 456 43 458 71
rect 466 43 468 71
rect 477 50 479 64
rect 487 50 489 64
rect 519 43 521 71
rect 529 43 531 71
rect 539 43 541 71
rect 557 43 559 68
rect 564 43 566 68
rect 574 46 576 59
rect 587 46 589 71
rect -203 -51 -201 -33
rect -176 -60 -174 -33
rect -166 -60 -164 -33
rect -159 -60 -157 -33
rect -149 -60 -147 -33
rect -139 -60 -137 -33
rect -114 -61 -112 -33
rect -104 -61 -102 -33
rect -94 -61 -92 -33
rect -84 -61 -82 -47
rect -74 -61 -72 -47
rect -54 -61 -52 -33
rect -44 -61 -42 -33
rect -34 -61 -32 -33
rect -23 -54 -21 -40
rect -13 -54 -11 -40
rect 17 -51 19 -33
rect 44 -60 46 -33
rect 54 -60 56 -33
rect 61 -60 63 -33
rect 71 -60 73 -33
rect 81 -60 83 -33
rect 106 -61 108 -33
rect 116 -61 118 -33
rect 126 -61 128 -33
rect 136 -61 138 -47
rect 146 -61 148 -47
rect 166 -61 168 -33
rect 176 -61 178 -33
rect 186 -61 188 -33
rect 197 -54 199 -40
rect 207 -54 209 -40
rect 234 -51 236 -33
rect 261 -60 263 -33
rect 271 -60 273 -33
rect 278 -60 280 -33
rect 288 -60 290 -33
rect 298 -60 300 -33
rect 323 -61 325 -33
rect 333 -61 335 -33
rect 343 -61 345 -33
rect 353 -61 355 -47
rect 363 -61 365 -47
rect 383 -61 385 -33
rect 393 -61 395 -33
rect 403 -61 405 -33
rect 414 -54 416 -40
rect 424 -54 426 -40
rect 462 -61 464 -33
rect 472 -61 474 -33
rect 482 -61 484 -33
rect 500 -58 502 -33
rect 507 -58 509 -33
rect 517 -49 519 -36
rect 530 -61 532 -36
<< polyct0 >>
rect 51 179 53 181
rect 91 179 93 181
rect 134 179 136 181
rect 238 179 240 181
rect 280 179 282 181
rect 324 179 326 181
rect 393 179 395 181
rect 437 179 439 181
rect 479 179 481 181
rect 520 179 522 181
rect 563 179 565 181
rect 603 179 605 181
rect 646 179 648 181
rect -66 116 -64 118
rect -24 116 -22 118
rect 22 116 24 118
rect 32 116 34 118
rect 88 123 90 125
rect 82 113 84 115
rect 204 116 206 118
rect 214 116 216 118
rect 254 116 256 118
rect 264 116 266 118
rect 274 116 276 118
rect 422 116 424 118
rect 432 116 434 118
rect 472 116 474 118
rect 482 116 484 118
rect 492 116 494 118
rect 560 116 562 118
rect 570 116 572 118
rect 626 123 628 125
rect 620 113 622 115
rect -183 36 -181 38
rect -50 36 -48 38
rect -40 36 -38 38
rect 0 36 2 38
rect 10 36 12 38
rect 20 36 22 38
rect 168 36 170 38
rect 178 36 180 38
rect 218 36 220 38
rect 228 36 230 38
rect 238 36 240 38
rect 388 36 390 38
rect 398 36 400 38
rect 438 36 440 38
rect 448 36 450 38
rect 458 36 460 38
rect 519 36 521 38
rect 529 36 531 38
rect 579 39 581 41
rect 585 29 587 31
rect -112 -28 -110 -26
rect -102 -28 -100 -26
rect -62 -28 -60 -26
rect -52 -28 -50 -26
rect -42 -28 -40 -26
rect 108 -28 110 -26
rect 118 -28 120 -26
rect 158 -28 160 -26
rect 168 -28 170 -26
rect 178 -28 180 -26
rect 325 -28 327 -26
rect 335 -28 337 -26
rect 375 -28 377 -26
rect 385 -28 387 -26
rect 395 -28 397 -26
rect 462 -28 464 -26
rect 472 -28 474 -26
rect 528 -21 530 -19
rect 522 -31 524 -29
<< polyct1 >>
rect 71 187 73 189
rect 61 179 63 181
rect 111 187 113 189
rect 101 179 103 181
rect 154 187 156 189
rect 144 179 146 181
rect 258 187 260 189
rect 248 179 250 181
rect 300 187 302 189
rect 290 179 292 181
rect 344 187 346 189
rect 334 179 336 181
rect 413 187 415 189
rect 403 179 405 181
rect 457 187 459 189
rect 447 179 449 181
rect 499 187 501 189
rect 489 179 491 181
rect 540 187 542 189
rect 530 179 532 181
rect 583 187 585 189
rect 573 179 575 181
rect 623 187 625 189
rect 613 179 615 181
rect 666 187 668 189
rect 656 179 658 181
rect -56 116 -54 118
rect -14 116 -12 118
rect -46 108 -44 110
rect 42 116 44 118
rect 49 116 51 118
rect 68 116 70 118
rect -4 108 -2 110
rect 115 116 117 118
rect 139 116 141 118
rect 165 116 167 118
rect 179 116 181 118
rect 244 122 246 124
rect 292 117 294 119
rect 240 102 242 104
rect 333 116 335 118
rect 357 116 359 118
rect 383 116 385 118
rect 397 116 399 118
rect 462 122 464 124
rect 510 117 512 119
rect 315 109 317 111
rect 458 102 460 104
rect 580 116 582 118
rect 587 116 589 118
rect 606 116 608 118
rect 533 109 535 111
rect -163 44 -161 46
rect -14 50 -12 52
rect -173 36 -171 38
rect -139 36 -137 38
rect -115 36 -113 38
rect -89 36 -87 38
rect -75 36 -73 38
rect 38 35 40 37
rect -10 30 -8 32
rect 61 43 63 45
rect 204 50 206 52
rect 79 36 81 38
rect 103 36 105 38
rect 129 36 131 38
rect 143 36 145 38
rect 256 35 258 37
rect 208 30 210 32
rect 279 43 281 45
rect 424 50 426 52
rect 299 36 301 38
rect 323 36 325 38
rect 349 36 351 38
rect 363 36 365 38
rect 476 35 478 37
rect 428 30 430 32
rect 499 43 501 45
rect 539 36 541 38
rect 546 36 548 38
rect 565 36 567 38
rect -201 -28 -199 -26
rect -177 -28 -175 -26
rect -151 -28 -149 -26
rect -137 -28 -135 -26
rect -72 -22 -70 -20
rect -24 -27 -22 -25
rect -76 -42 -74 -40
rect 19 -28 21 -26
rect 43 -28 45 -26
rect 69 -28 71 -26
rect 83 -28 85 -26
rect 148 -22 150 -20
rect 196 -27 198 -25
rect -1 -35 1 -33
rect 144 -42 146 -40
rect 236 -28 238 -26
rect 260 -28 262 -26
rect 286 -28 288 -26
rect 300 -28 302 -26
rect 365 -22 367 -20
rect 413 -27 415 -25
rect 219 -35 221 -33
rect 361 -42 363 -40
rect 482 -28 484 -26
rect 489 -28 491 -26
rect 508 -28 510 -26
rect 436 -35 438 -33
<< ndifct0 >>
rect 74 163 76 165
rect 114 163 116 165
rect 157 163 159 165
rect 261 163 263 165
rect 303 163 305 165
rect 347 163 349 165
rect 416 163 418 165
rect 460 163 462 165
rect 502 163 504 165
rect 543 163 545 165
rect 586 163 588 165
rect 626 163 628 165
rect 669 163 671 165
rect -43 132 -41 134
rect -1 132 1 134
rect 28 139 30 141
rect 45 132 47 134
rect 55 132 57 134
rect 55 125 57 127
rect 65 125 67 127
rect 75 133 77 135
rect 85 136 87 138
rect 132 133 134 135
rect 122 128 124 130
rect 171 131 173 133
rect 181 131 183 133
rect 236 139 238 141
rect 225 131 227 133
rect 247 131 249 133
rect 277 132 279 134
rect 287 131 289 133
rect 297 133 299 135
rect 350 133 352 135
rect 308 125 310 127
rect 340 128 342 130
rect 389 131 391 133
rect 399 131 401 133
rect 454 139 456 141
rect 443 131 445 133
rect 465 131 467 133
rect 495 132 497 134
rect 505 131 507 133
rect 515 133 517 135
rect 566 139 568 141
rect 526 125 528 127
rect 583 132 585 134
rect 593 132 595 134
rect 593 125 595 127
rect 603 125 605 127
rect 613 133 615 135
rect 623 136 625 138
rect -132 24 -130 26
rect -160 20 -158 22
rect -122 19 -120 21
rect -83 21 -81 23
rect -73 21 -71 23
rect -29 21 -27 23
rect -18 13 -16 15
rect -7 21 -5 23
rect 23 20 25 22
rect 33 21 35 23
rect 43 19 45 21
rect 54 27 56 29
rect 86 24 88 26
rect 96 19 98 21
rect 135 21 137 23
rect 145 21 147 23
rect 189 21 191 23
rect 200 13 202 15
rect 211 21 213 23
rect 241 20 243 22
rect 251 21 253 23
rect 261 19 263 21
rect 272 27 274 29
rect 306 24 308 26
rect 316 19 318 21
rect 355 21 357 23
rect 365 21 367 23
rect 409 21 411 23
rect 420 13 422 15
rect 431 21 433 23
rect 461 20 463 22
rect 471 21 473 23
rect 481 19 483 21
rect 492 27 494 29
rect 525 13 527 15
rect 552 27 554 29
rect 542 20 544 22
rect 552 20 554 22
rect 562 27 564 29
rect 572 19 574 21
rect 582 16 584 18
rect -184 -11 -182 -9
rect -194 -16 -192 -14
rect -145 -13 -143 -11
rect -135 -13 -133 -11
rect -80 -5 -78 -3
rect -91 -13 -89 -11
rect -69 -13 -67 -11
rect -39 -12 -37 -10
rect -29 -13 -27 -11
rect -19 -11 -17 -9
rect 36 -11 38 -9
rect -8 -19 -6 -17
rect 26 -16 28 -14
rect 75 -13 77 -11
rect 85 -13 87 -11
rect 140 -5 142 -3
rect 129 -13 131 -11
rect 151 -13 153 -11
rect 181 -12 183 -10
rect 191 -13 193 -11
rect 201 -11 203 -9
rect 253 -11 255 -9
rect 212 -19 214 -17
rect 243 -16 245 -14
rect 292 -13 294 -11
rect 302 -13 304 -11
rect 357 -5 359 -3
rect 346 -13 348 -11
rect 368 -13 370 -11
rect 398 -12 400 -10
rect 408 -13 410 -11
rect 418 -11 420 -9
rect 468 -5 470 -3
rect 429 -19 431 -17
rect 485 -12 487 -10
rect 495 -12 497 -10
rect 495 -19 497 -17
rect 505 -19 507 -17
rect 515 -11 517 -9
rect 525 -8 527 -6
<< ndifct1 >>
rect 44 165 46 167
rect 84 165 86 167
rect 127 165 129 167
rect 55 153 57 155
rect 231 165 233 167
rect 95 153 97 155
rect 273 165 275 167
rect 138 153 140 155
rect 317 165 319 167
rect 242 153 244 155
rect 386 165 388 167
rect 284 153 286 155
rect 430 165 432 167
rect 328 153 330 155
rect 472 165 474 167
rect 397 153 399 155
rect 513 165 515 167
rect 441 153 443 155
rect 556 165 558 167
rect 483 153 485 155
rect 596 165 598 167
rect 524 153 526 155
rect 639 165 641 167
rect 567 153 569 155
rect 607 153 609 155
rect 650 153 652 155
rect -62 142 -60 144
rect -20 142 -18 144
rect -73 130 -71 132
rect -31 130 -29 132
rect 17 132 19 134
rect 143 142 145 144
rect 95 132 97 134
rect 108 125 110 127
rect 197 142 199 144
rect 161 125 163 127
rect 215 132 217 134
rect 259 142 261 144
rect 361 142 363 144
rect 326 125 328 127
rect 415 142 417 144
rect 379 125 381 127
rect 433 132 435 134
rect 477 142 479 144
rect 555 132 557 134
rect 633 132 635 134
rect -190 22 -188 24
rect -146 27 -144 29
rect -93 27 -91 29
rect -179 10 -177 12
rect -111 10 -109 12
rect -39 20 -37 22
rect -57 10 -55 12
rect 72 27 74 29
rect 5 10 7 12
rect 125 27 127 29
rect 107 10 109 12
rect 179 20 181 22
rect 161 10 163 12
rect 292 27 294 29
rect 223 10 225 12
rect 345 27 347 29
rect 327 10 329 12
rect 399 20 401 22
rect 381 10 383 12
rect 514 20 516 22
rect 443 10 445 12
rect 592 20 594 22
rect -173 -2 -171 0
rect -208 -19 -206 -17
rect -119 -2 -117 0
rect -155 -19 -153 -17
rect -101 -12 -99 -10
rect -57 -2 -55 0
rect 47 -2 49 0
rect 12 -19 14 -17
rect 101 -2 103 0
rect 65 -19 67 -17
rect 119 -12 121 -10
rect 163 -2 165 0
rect 264 -2 266 0
rect 229 -19 231 -17
rect 318 -2 320 0
rect 282 -19 284 -17
rect 336 -12 338 -10
rect 380 -2 382 0
rect 457 -12 459 -10
rect 535 -12 537 -10
<< ntiect1 >>
rect 45 213 47 215
rect 85 213 87 215
rect 128 213 130 215
rect 232 213 234 215
rect 274 213 276 215
rect 318 213 320 215
rect 387 213 389 215
rect 431 213 433 215
rect 473 213 475 215
rect 514 213 516 215
rect 557 213 559 215
rect 597 213 599 215
rect 640 213 642 215
rect -72 82 -70 84
rect -30 82 -28 84
rect 109 82 111 84
rect 121 82 123 84
rect 314 82 316 84
rect 327 82 329 84
rect 339 82 341 84
rect 532 82 534 84
rect -189 70 -187 72
rect -145 70 -143 72
rect -133 70 -131 72
rect 60 70 62 72
rect 73 70 75 72
rect 85 70 87 72
rect 278 70 280 72
rect 293 70 295 72
rect 305 70 307 72
rect 498 70 500 72
rect -207 -62 -205 -60
rect -195 -62 -193 -60
rect -2 -62 0 -60
rect 13 -62 15 -60
rect 25 -62 27 -60
rect 218 -62 220 -60
rect 230 -62 232 -60
rect 242 -62 244 -60
rect 435 -62 437 -60
<< ptiect1 >>
rect 45 153 47 155
rect 85 153 87 155
rect 128 153 130 155
rect 232 153 234 155
rect 274 153 276 155
rect 318 153 320 155
rect 387 153 389 155
rect 431 153 433 155
rect 473 153 475 155
rect 514 153 516 155
rect 557 153 559 155
rect 597 153 599 155
rect 640 153 642 155
rect -72 142 -70 144
rect -30 142 -28 144
rect 109 142 111 144
rect 121 142 123 144
rect 314 142 316 144
rect 327 142 329 144
rect 339 142 341 144
rect 532 142 534 144
rect -189 10 -187 12
rect -145 10 -143 12
rect -133 10 -131 12
rect 60 10 62 12
rect 73 10 75 12
rect 85 10 87 12
rect 278 10 280 12
rect 293 10 295 12
rect 305 10 307 12
rect 498 10 500 12
rect -207 -2 -205 0
rect -195 -2 -193 0
rect -2 -2 0 0
rect 13 -2 15 0
rect 25 -2 27 0
rect 218 -2 220 0
rect 230 -2 232 0
rect 242 -2 244 0
rect 435 -2 437 0
<< pdifct0 >>
rect 54 201 56 203
rect 64 203 66 205
rect 64 196 66 198
rect 74 203 76 205
rect 94 201 96 203
rect 104 203 106 205
rect 104 196 106 198
rect 114 203 116 205
rect 137 201 139 203
rect 147 203 149 205
rect 147 196 149 198
rect 157 203 159 205
rect 241 201 243 203
rect 251 203 253 205
rect 251 196 253 198
rect 261 203 263 205
rect 283 201 285 203
rect 293 203 295 205
rect 293 196 295 198
rect 303 203 305 205
rect 327 201 329 203
rect 337 203 339 205
rect 337 196 339 198
rect 347 203 349 205
rect 396 201 398 203
rect 406 203 408 205
rect 406 196 408 198
rect 416 203 418 205
rect 440 201 442 203
rect 450 203 452 205
rect 450 196 452 198
rect 460 203 462 205
rect 482 201 484 203
rect 492 203 494 205
rect 492 196 494 198
rect 502 203 504 205
rect 523 201 525 203
rect 533 203 535 205
rect 533 196 535 198
rect 543 203 545 205
rect 566 201 568 203
rect 576 203 578 205
rect 576 196 578 198
rect 586 203 588 205
rect 606 201 608 203
rect 616 203 618 205
rect 616 196 618 198
rect 626 203 628 205
rect 649 201 651 203
rect 659 203 661 205
rect 659 196 661 198
rect 669 203 671 205
rect -63 94 -61 96
rect -53 99 -51 101
rect -53 92 -51 94
rect -43 92 -41 94
rect -21 94 -19 96
rect -11 99 -9 101
rect -11 92 -9 94
rect -1 92 1 94
rect 27 92 29 94
rect 27 85 29 87
rect 37 100 39 102
rect 37 93 39 95
rect 49 92 51 94
rect 49 85 51 87
rect 72 104 74 106
rect 84 85 86 87
rect 119 92 121 94
rect 135 99 137 101
rect 135 92 137 94
rect 145 93 147 95
rect 145 86 147 88
rect 172 91 174 93
rect 182 94 184 96
rect 197 92 199 94
rect 182 86 184 88
rect 217 107 219 109
rect 217 100 219 102
rect 227 85 229 87
rect 237 92 239 94
rect 247 92 249 94
rect 257 92 259 94
rect 247 85 249 87
rect 267 100 269 102
rect 277 107 279 109
rect 277 100 279 102
rect 298 100 300 102
rect 308 92 310 94
rect 287 85 289 87
rect 337 92 339 94
rect 353 99 355 101
rect 353 92 355 94
rect 363 93 365 95
rect 363 86 365 88
rect 390 91 392 93
rect 400 94 402 96
rect 415 92 417 94
rect 400 86 402 88
rect 435 107 437 109
rect 435 100 437 102
rect 445 85 447 87
rect 455 92 457 94
rect 465 92 467 94
rect 475 92 477 94
rect 465 85 467 87
rect 485 100 487 102
rect 495 107 497 109
rect 495 100 497 102
rect 516 100 518 102
rect 526 92 528 94
rect 505 85 507 87
rect 565 92 567 94
rect 565 85 567 87
rect 575 100 577 102
rect 575 93 577 95
rect 587 92 589 94
rect 587 85 589 87
rect 610 104 612 106
rect 622 85 624 87
rect -180 58 -178 60
rect -170 60 -168 62
rect -170 53 -168 55
rect -160 60 -158 62
rect -135 60 -133 62
rect -119 60 -117 62
rect -119 53 -117 55
rect -109 66 -107 68
rect -109 59 -107 61
rect -82 61 -80 63
rect -72 66 -70 68
rect -72 58 -70 60
rect -57 60 -55 62
rect -37 52 -35 54
rect -37 45 -35 47
rect -27 67 -25 69
rect -17 60 -15 62
rect -7 67 -5 69
rect -7 60 -5 62
rect 3 60 5 62
rect 13 52 15 54
rect 23 52 25 54
rect 23 45 25 47
rect 33 67 35 69
rect 44 52 46 54
rect 54 60 56 62
rect 83 60 85 62
rect 99 60 101 62
rect 99 53 101 55
rect 109 66 111 68
rect 109 59 111 61
rect 136 61 138 63
rect 146 66 148 68
rect 146 58 148 60
rect 161 60 163 62
rect 181 52 183 54
rect 181 45 183 47
rect 191 67 193 69
rect 201 60 203 62
rect 211 67 213 69
rect 211 60 213 62
rect 221 60 223 62
rect 231 52 233 54
rect 241 52 243 54
rect 241 45 243 47
rect 251 67 253 69
rect 262 52 264 54
rect 272 60 274 62
rect 303 60 305 62
rect 319 60 321 62
rect 319 53 321 55
rect 329 66 331 68
rect 329 59 331 61
rect 356 61 358 63
rect 366 66 368 68
rect 366 58 368 60
rect 381 60 383 62
rect 401 52 403 54
rect 401 45 403 47
rect 411 67 413 69
rect 421 60 423 62
rect 431 67 433 69
rect 431 60 433 62
rect 441 60 443 62
rect 451 52 453 54
rect 461 52 463 54
rect 461 45 463 47
rect 471 67 473 69
rect 482 52 484 54
rect 492 60 494 62
rect 524 67 526 69
rect 524 60 526 62
rect 534 59 536 61
rect 534 52 536 54
rect 546 67 548 69
rect 546 60 548 62
rect 581 67 583 69
rect 569 48 571 50
rect -197 -52 -195 -50
rect -181 -45 -179 -43
rect -181 -52 -179 -50
rect -171 -51 -169 -49
rect -171 -58 -169 -56
rect -144 -53 -142 -51
rect -134 -50 -132 -48
rect -119 -52 -117 -50
rect -134 -58 -132 -56
rect -99 -37 -97 -35
rect -99 -44 -97 -42
rect -89 -59 -87 -57
rect -79 -52 -77 -50
rect -69 -52 -67 -50
rect -59 -52 -57 -50
rect -69 -59 -67 -57
rect -49 -44 -47 -42
rect -39 -37 -37 -35
rect -39 -44 -37 -42
rect -18 -44 -16 -42
rect -8 -52 -6 -50
rect -29 -59 -27 -57
rect 23 -52 25 -50
rect 39 -45 41 -43
rect 39 -52 41 -50
rect 49 -51 51 -49
rect 49 -58 51 -56
rect 76 -53 78 -51
rect 86 -50 88 -48
rect 101 -52 103 -50
rect 86 -58 88 -56
rect 121 -37 123 -35
rect 121 -44 123 -42
rect 131 -59 133 -57
rect 141 -52 143 -50
rect 151 -52 153 -50
rect 161 -52 163 -50
rect 151 -59 153 -57
rect 171 -44 173 -42
rect 181 -37 183 -35
rect 181 -44 183 -42
rect 202 -44 204 -42
rect 212 -52 214 -50
rect 191 -59 193 -57
rect 240 -52 242 -50
rect 256 -45 258 -43
rect 256 -52 258 -50
rect 266 -51 268 -49
rect 266 -58 268 -56
rect 293 -53 295 -51
rect 303 -50 305 -48
rect 318 -52 320 -50
rect 303 -58 305 -56
rect 338 -37 340 -35
rect 338 -44 340 -42
rect 348 -59 350 -57
rect 358 -52 360 -50
rect 368 -52 370 -50
rect 378 -52 380 -50
rect 368 -59 370 -57
rect 388 -44 390 -42
rect 398 -37 400 -35
rect 398 -44 400 -42
rect 419 -44 421 -42
rect 429 -52 431 -50
rect 408 -59 410 -57
rect 467 -52 469 -50
rect 467 -59 469 -57
rect 477 -44 479 -42
rect 477 -51 479 -49
rect 489 -52 491 -50
rect 489 -59 491 -57
rect 512 -40 514 -38
rect 524 -59 526 -57
<< pdifct1 >>
rect 44 196 46 198
rect 44 189 46 191
rect 84 196 86 198
rect 84 189 86 191
rect 127 196 129 198
rect 127 189 129 191
rect 231 196 233 198
rect 231 189 233 191
rect 273 196 275 198
rect 273 189 275 191
rect 317 196 319 198
rect 317 189 319 191
rect 386 196 388 198
rect 386 189 388 191
rect 430 196 432 198
rect 430 189 432 191
rect 472 196 474 198
rect 472 189 474 191
rect 513 196 515 198
rect 513 189 515 191
rect 556 196 558 198
rect 556 189 558 191
rect 596 196 598 198
rect 596 189 598 191
rect 639 196 641 198
rect 639 189 641 191
rect -73 106 -71 108
rect -73 99 -71 101
rect -31 106 -29 108
rect -31 99 -29 101
rect 17 107 19 109
rect 17 100 19 102
rect 95 104 97 106
rect 95 97 97 99
rect 108 107 110 109
rect 108 100 110 102
rect 162 107 164 109
rect 162 100 164 102
rect 207 100 209 102
rect 326 107 328 109
rect 326 100 328 102
rect 380 107 382 109
rect 380 100 382 102
rect 425 100 427 102
rect 555 107 557 109
rect 555 100 557 102
rect 633 104 635 106
rect 633 97 635 99
rect -190 53 -188 55
rect -190 46 -188 48
rect -146 52 -144 54
rect -146 45 -144 47
rect -92 52 -90 54
rect -92 45 -90 47
rect -47 52 -45 54
rect 72 52 74 54
rect 72 45 74 47
rect 126 52 128 54
rect 126 45 128 47
rect 171 52 173 54
rect 292 52 294 54
rect 292 45 294 47
rect 346 52 348 54
rect 346 45 348 47
rect 391 52 393 54
rect 514 52 516 54
rect 514 45 516 47
rect 592 55 594 57
rect 592 48 594 50
rect -208 -37 -206 -35
rect -208 -44 -206 -42
rect -154 -37 -152 -35
rect -154 -44 -152 -42
rect -109 -44 -107 -42
rect 12 -37 14 -35
rect 12 -44 14 -42
rect 66 -37 68 -35
rect 66 -44 68 -42
rect 111 -44 113 -42
rect 229 -37 231 -35
rect 229 -44 231 -42
rect 283 -37 285 -35
rect 283 -44 285 -42
rect 328 -44 330 -42
rect 457 -37 459 -35
rect 457 -44 459 -42
rect 535 -40 537 -38
rect 535 -47 537 -45
<< alu0 >>
rect 52 203 58 212
rect 52 201 54 203
rect 56 201 58 203
rect 52 200 58 201
rect 63 205 67 207
rect 63 203 64 205
rect 66 203 67 205
rect 63 198 67 203
rect 72 205 78 212
rect 72 203 74 205
rect 76 203 78 205
rect 72 202 78 203
rect 92 203 98 212
rect 92 201 94 203
rect 96 201 98 203
rect 92 200 98 201
rect 103 205 107 207
rect 103 203 104 205
rect 106 203 107 205
rect 63 197 64 198
rect 50 196 64 197
rect 66 196 67 198
rect 50 193 67 196
rect 50 181 54 193
rect 103 198 107 203
rect 112 205 118 212
rect 112 203 114 205
rect 116 203 118 205
rect 112 202 118 203
rect 135 203 141 212
rect 135 201 137 203
rect 139 201 141 203
rect 135 200 141 201
rect 146 205 150 207
rect 146 203 147 205
rect 149 203 150 205
rect 103 197 104 198
rect 90 196 104 197
rect 106 196 107 198
rect 90 193 107 196
rect 50 179 51 181
rect 53 179 54 181
rect 50 174 54 179
rect 50 170 62 174
rect 46 167 47 169
rect 58 166 62 170
rect 90 181 94 193
rect 146 198 150 203
rect 155 205 161 212
rect 155 203 157 205
rect 159 203 161 205
rect 155 202 161 203
rect 239 203 245 212
rect 239 201 241 203
rect 243 201 245 203
rect 239 200 245 201
rect 250 205 254 207
rect 250 203 251 205
rect 253 203 254 205
rect 146 197 147 198
rect 133 196 147 197
rect 149 196 150 198
rect 133 193 150 196
rect 90 179 91 181
rect 93 179 94 181
rect 90 174 94 179
rect 90 170 102 174
rect 86 167 87 169
rect 58 165 78 166
rect 58 163 74 165
rect 76 163 78 165
rect 58 162 78 163
rect 98 166 102 170
rect 133 181 137 193
rect 250 198 254 203
rect 259 205 265 212
rect 259 203 261 205
rect 263 203 265 205
rect 259 202 265 203
rect 281 203 287 212
rect 281 201 283 203
rect 285 201 287 203
rect 281 200 287 201
rect 292 205 296 207
rect 292 203 293 205
rect 295 203 296 205
rect 250 197 251 198
rect 237 196 251 197
rect 253 196 254 198
rect 237 193 254 196
rect 133 179 134 181
rect 136 179 137 181
rect 133 174 137 179
rect 133 170 145 174
rect 129 167 130 169
rect 98 165 118 166
rect 98 163 114 165
rect 116 163 118 165
rect 98 162 118 163
rect 141 166 145 170
rect 237 181 241 193
rect 292 198 296 203
rect 301 205 307 212
rect 301 203 303 205
rect 305 203 307 205
rect 301 202 307 203
rect 325 203 331 212
rect 325 201 327 203
rect 329 201 331 203
rect 325 200 331 201
rect 336 205 340 207
rect 336 203 337 205
rect 339 203 340 205
rect 292 197 293 198
rect 279 196 293 197
rect 295 196 296 198
rect 279 193 296 196
rect 237 179 238 181
rect 240 179 241 181
rect 237 174 241 179
rect 237 170 249 174
rect 233 167 234 169
rect 141 165 161 166
rect 141 163 157 165
rect 159 163 161 165
rect 141 162 161 163
rect 245 166 249 170
rect 279 181 283 193
rect 336 198 340 203
rect 345 205 351 212
rect 345 203 347 205
rect 349 203 351 205
rect 345 202 351 203
rect 394 203 400 212
rect 394 201 396 203
rect 398 201 400 203
rect 394 200 400 201
rect 405 205 409 207
rect 405 203 406 205
rect 408 203 409 205
rect 336 197 337 198
rect 323 196 337 197
rect 339 196 340 198
rect 323 193 340 196
rect 279 179 280 181
rect 282 179 283 181
rect 279 174 283 179
rect 279 170 291 174
rect 275 167 276 169
rect 245 165 265 166
rect 245 163 261 165
rect 263 163 265 165
rect 245 162 265 163
rect 287 166 291 170
rect 323 181 327 193
rect 405 198 409 203
rect 414 205 420 212
rect 414 203 416 205
rect 418 203 420 205
rect 414 202 420 203
rect 438 203 444 212
rect 438 201 440 203
rect 442 201 444 203
rect 438 200 444 201
rect 449 205 453 207
rect 449 203 450 205
rect 452 203 453 205
rect 405 197 406 198
rect 392 196 406 197
rect 408 196 409 198
rect 392 193 409 196
rect 323 179 324 181
rect 326 179 327 181
rect 323 174 327 179
rect 323 170 335 174
rect 319 167 320 169
rect 287 165 307 166
rect 287 163 303 165
rect 305 163 307 165
rect 287 162 307 163
rect 331 166 335 170
rect 392 181 396 193
rect 449 198 453 203
rect 458 205 464 212
rect 458 203 460 205
rect 462 203 464 205
rect 458 202 464 203
rect 480 203 486 212
rect 480 201 482 203
rect 484 201 486 203
rect 480 200 486 201
rect 491 205 495 207
rect 491 203 492 205
rect 494 203 495 205
rect 449 197 450 198
rect 436 196 450 197
rect 452 196 453 198
rect 436 193 453 196
rect 392 179 393 181
rect 395 179 396 181
rect 392 174 396 179
rect 392 170 404 174
rect 388 167 389 169
rect 331 165 351 166
rect 331 163 347 165
rect 349 163 351 165
rect 331 162 351 163
rect 400 166 404 170
rect 436 181 440 193
rect 491 198 495 203
rect 500 205 506 212
rect 500 203 502 205
rect 504 203 506 205
rect 500 202 506 203
rect 521 203 527 212
rect 521 201 523 203
rect 525 201 527 203
rect 521 200 527 201
rect 532 205 536 207
rect 532 203 533 205
rect 535 203 536 205
rect 491 197 492 198
rect 478 196 492 197
rect 494 196 495 198
rect 478 193 495 196
rect 436 179 437 181
rect 439 179 440 181
rect 436 174 440 179
rect 436 170 448 174
rect 432 167 433 169
rect 400 165 420 166
rect 400 163 416 165
rect 418 163 420 165
rect 400 162 420 163
rect 444 166 448 170
rect 478 181 482 193
rect 532 198 536 203
rect 541 205 547 212
rect 541 203 543 205
rect 545 203 547 205
rect 541 202 547 203
rect 564 203 570 212
rect 564 201 566 203
rect 568 201 570 203
rect 564 200 570 201
rect 575 205 579 207
rect 575 203 576 205
rect 578 203 579 205
rect 532 197 533 198
rect 519 196 533 197
rect 535 196 536 198
rect 519 193 536 196
rect 478 179 479 181
rect 481 179 482 181
rect 478 174 482 179
rect 478 170 490 174
rect 474 167 475 169
rect 444 165 464 166
rect 444 163 460 165
rect 462 163 464 165
rect 444 162 464 163
rect 486 166 490 170
rect 519 181 523 193
rect 575 198 579 203
rect 584 205 590 212
rect 584 203 586 205
rect 588 203 590 205
rect 584 202 590 203
rect 604 203 610 212
rect 604 201 606 203
rect 608 201 610 203
rect 604 200 610 201
rect 615 205 619 207
rect 615 203 616 205
rect 618 203 619 205
rect 575 197 576 198
rect 562 196 576 197
rect 578 196 579 198
rect 562 193 579 196
rect 519 179 520 181
rect 522 179 523 181
rect 519 174 523 179
rect 519 170 531 174
rect 515 167 516 169
rect 486 165 506 166
rect 486 163 502 165
rect 504 163 506 165
rect 486 162 506 163
rect 527 166 531 170
rect 562 181 566 193
rect 615 198 619 203
rect 624 205 630 212
rect 624 203 626 205
rect 628 203 630 205
rect 624 202 630 203
rect 647 203 653 212
rect 647 201 649 203
rect 651 201 653 203
rect 647 200 653 201
rect 658 205 662 207
rect 658 203 659 205
rect 661 203 662 205
rect 615 197 616 198
rect 602 196 616 197
rect 618 196 619 198
rect 602 193 619 196
rect 562 179 563 181
rect 565 179 566 181
rect 562 174 566 179
rect 562 170 574 174
rect 558 167 559 169
rect 527 165 547 166
rect 527 163 543 165
rect 545 163 547 165
rect 527 162 547 163
rect 570 166 574 170
rect 602 181 606 193
rect 658 198 662 203
rect 667 205 673 212
rect 667 203 669 205
rect 671 203 673 205
rect 667 202 673 203
rect 658 197 659 198
rect 645 196 659 197
rect 661 196 662 198
rect 645 193 662 196
rect 602 179 603 181
rect 605 179 606 181
rect 602 174 606 179
rect 602 170 614 174
rect 598 167 599 169
rect 570 165 590 166
rect 570 163 586 165
rect 588 163 590 165
rect 570 162 590 163
rect 610 166 614 170
rect 645 181 649 193
rect 645 179 646 181
rect 648 179 649 181
rect 645 174 649 179
rect 645 170 657 174
rect 641 167 642 169
rect 610 165 630 166
rect 610 163 626 165
rect 628 163 630 165
rect 610 162 630 163
rect 653 166 657 170
rect 653 165 673 166
rect 653 163 669 165
rect 671 163 673 165
rect 653 162 673 163
rect 26 139 28 141
rect 30 139 32 141
rect 26 138 32 139
rect 84 138 88 141
rect 84 136 85 138
rect 87 136 88 138
rect -59 134 -39 135
rect -59 132 -43 134
rect -41 132 -39 134
rect -59 131 -39 132
rect 54 135 79 136
rect -71 128 -70 130
rect -59 127 -55 131
rect -17 134 3 135
rect -17 132 -1 134
rect 1 132 3 134
rect -17 131 3 132
rect 39 134 49 135
rect 39 132 45 134
rect 47 132 49 134
rect 39 131 49 132
rect 54 134 75 135
rect 54 132 55 134
rect 57 133 75 134
rect 77 133 79 135
rect 84 134 88 136
rect 57 132 79 133
rect -67 123 -55 127
rect -67 118 -63 123
rect -67 116 -66 118
rect -64 116 -63 118
rect -67 104 -63 116
rect -67 101 -50 104
rect -67 100 -53 101
rect -54 99 -53 100
rect -51 99 -50 101
rect -65 96 -59 97
rect -65 94 -63 96
rect -61 94 -59 96
rect -65 85 -59 94
rect -54 94 -50 99
rect -29 128 -28 130
rect -17 127 -13 131
rect -25 123 -13 127
rect -25 118 -21 123
rect -25 116 -24 118
rect -22 116 -21 118
rect -25 104 -21 116
rect 39 127 43 131
rect 23 123 43 127
rect 23 120 27 123
rect 21 118 27 120
rect 21 116 22 118
rect 24 116 27 118
rect 21 114 27 116
rect -25 101 -8 104
rect -25 100 -11 101
rect -12 99 -11 100
rect -9 99 -8 101
rect -23 96 -17 97
rect -54 92 -53 94
rect -51 92 -50 94
rect -54 90 -50 92
rect -45 94 -39 95
rect -45 92 -43 94
rect -41 92 -39 94
rect -45 85 -39 92
rect -23 94 -21 96
rect -19 94 -17 96
rect -23 85 -17 94
rect -12 94 -8 99
rect 23 103 27 114
rect 31 118 35 120
rect 54 127 58 132
rect 54 125 55 127
rect 57 125 58 127
rect 54 123 58 125
rect 63 127 78 128
rect 63 125 65 127
rect 67 126 78 127
rect 67 125 92 126
rect 63 124 88 125
rect 74 123 88 124
rect 90 123 92 125
rect 74 122 92 123
rect 31 116 32 118
rect 34 116 35 118
rect 31 111 35 116
rect 74 111 78 122
rect 71 107 78 111
rect 81 115 85 117
rect 81 113 82 115
rect 84 113 85 115
rect 71 106 75 107
rect 71 104 72 106
rect 74 104 75 106
rect 23 102 63 103
rect 71 102 75 104
rect 81 103 85 113
rect 23 100 37 102
rect 39 100 63 102
rect 23 99 63 100
rect 79 99 85 103
rect 36 95 40 99
rect 59 95 83 99
rect 121 130 125 141
rect 130 135 175 136
rect 130 133 132 135
rect 134 133 175 135
rect 130 132 171 133
rect 169 131 171 132
rect 173 131 175 133
rect 169 130 175 131
rect 179 133 185 141
rect 234 139 236 141
rect 238 139 240 141
rect 234 138 240 139
rect 296 135 300 141
rect 179 131 181 133
rect 183 131 185 133
rect 179 130 185 131
rect 224 133 228 135
rect 255 134 281 135
rect 224 131 225 133
rect 227 131 228 133
rect 110 123 111 129
rect 121 128 122 130
rect 124 128 125 130
rect 121 126 125 128
rect 110 104 111 111
rect 134 101 156 103
rect 134 99 135 101
rect 137 99 156 101
rect -12 92 -11 94
rect -9 92 -8 94
rect -12 90 -8 92
rect -3 94 3 95
rect -3 92 -1 94
rect 1 92 3 94
rect -3 85 3 92
rect 25 94 31 95
rect 25 92 27 94
rect 29 92 31 94
rect 25 87 31 92
rect 36 93 37 95
rect 39 93 40 95
rect 36 91 40 93
rect 47 94 53 95
rect 47 92 49 94
rect 51 92 53 94
rect 25 85 27 87
rect 29 85 31 87
rect 47 87 53 92
rect 117 94 123 95
rect 117 92 119 94
rect 121 92 123 94
rect 47 85 49 87
rect 51 85 53 87
rect 82 87 88 88
rect 82 85 84 87
rect 86 85 88 87
rect 117 85 123 92
rect 134 94 138 99
rect 134 92 135 94
rect 137 92 138 94
rect 134 90 138 92
rect 143 95 149 96
rect 143 93 145 95
rect 147 93 149 95
rect 143 88 149 93
rect 152 94 156 99
rect 224 127 228 131
rect 203 123 228 127
rect 234 133 251 134
rect 234 131 247 133
rect 249 131 251 133
rect 234 130 251 131
rect 255 132 277 134
rect 279 132 281 134
rect 255 131 281 132
rect 286 133 290 135
rect 286 131 287 133
rect 289 131 290 133
rect 296 133 297 135
rect 299 133 300 135
rect 296 131 300 133
rect 203 118 207 123
rect 234 119 238 130
rect 203 116 204 118
rect 206 116 207 118
rect 203 110 207 116
rect 212 118 238 119
rect 212 116 214 118
rect 216 116 238 118
rect 212 115 238 116
rect 255 119 259 131
rect 286 127 290 131
rect 307 127 311 129
rect 203 109 221 110
rect 203 107 217 109
rect 219 107 221 109
rect 203 106 221 107
rect 215 102 221 106
rect 215 100 217 102
rect 219 100 221 102
rect 215 99 221 100
rect 181 96 185 98
rect 181 94 182 96
rect 184 94 185 96
rect 225 95 229 115
rect 252 118 259 119
rect 252 116 254 118
rect 256 116 259 118
rect 252 115 259 116
rect 255 103 259 115
rect 263 123 290 127
rect 263 118 267 123
rect 263 116 264 118
rect 266 116 267 118
rect 263 111 267 116
rect 272 118 287 119
rect 272 116 274 118
rect 276 116 287 118
rect 272 115 287 116
rect 263 109 280 111
rect 263 107 277 109
rect 279 107 280 109
rect 255 102 271 103
rect 255 100 267 102
rect 269 100 271 102
rect 255 99 271 100
rect 276 102 280 107
rect 276 100 277 102
rect 279 100 280 102
rect 276 98 280 100
rect 283 102 287 115
rect 307 125 308 127
rect 310 125 311 127
rect 307 111 311 125
rect 339 130 343 141
rect 348 135 393 136
rect 348 133 350 135
rect 352 133 393 135
rect 348 132 389 133
rect 387 131 389 132
rect 391 131 393 133
rect 387 130 393 131
rect 397 133 403 141
rect 452 139 454 141
rect 456 139 458 141
rect 452 138 458 139
rect 514 135 518 141
rect 564 139 566 141
rect 568 139 570 141
rect 564 138 570 139
rect 622 138 626 141
rect 622 136 623 138
rect 625 136 626 138
rect 592 135 617 136
rect 397 131 399 133
rect 401 131 403 133
rect 397 130 403 131
rect 442 133 446 135
rect 473 134 499 135
rect 442 131 443 133
rect 445 131 446 133
rect 297 107 311 111
rect 297 102 301 107
rect 283 100 298 102
rect 300 100 301 102
rect 283 98 301 100
rect 328 123 329 129
rect 339 128 340 130
rect 342 128 343 130
rect 339 126 343 128
rect 328 104 329 111
rect 352 101 374 103
rect 352 99 353 101
rect 355 99 374 101
rect 283 95 287 98
rect 152 93 176 94
rect 152 91 172 93
rect 174 91 176 93
rect 152 90 176 91
rect 143 86 145 88
rect 147 86 149 88
rect 143 85 149 86
rect 181 88 185 94
rect 195 94 241 95
rect 195 92 197 94
rect 199 92 237 94
rect 239 92 241 94
rect 195 91 241 92
rect 245 94 251 95
rect 245 92 247 94
rect 249 92 251 94
rect 181 86 182 88
rect 184 86 185 88
rect 181 85 185 86
rect 225 87 231 88
rect 225 85 227 87
rect 229 85 231 87
rect 245 87 251 92
rect 255 94 287 95
rect 255 92 257 94
rect 259 92 287 94
rect 255 91 287 92
rect 306 94 312 95
rect 306 92 308 94
rect 310 92 312 94
rect 245 85 247 87
rect 249 85 251 87
rect 285 87 291 88
rect 285 85 287 87
rect 289 85 291 87
rect 306 85 312 92
rect 335 94 341 95
rect 335 92 337 94
rect 339 92 341 94
rect 335 85 341 92
rect 352 94 356 99
rect 352 92 353 94
rect 355 92 356 94
rect 352 90 356 92
rect 361 95 367 96
rect 361 93 363 95
rect 365 93 367 95
rect 361 88 367 93
rect 370 94 374 99
rect 442 127 446 131
rect 421 123 446 127
rect 452 133 469 134
rect 452 131 465 133
rect 467 131 469 133
rect 452 130 469 131
rect 473 132 495 134
rect 497 132 499 134
rect 473 131 499 132
rect 504 133 508 135
rect 504 131 505 133
rect 507 131 508 133
rect 514 133 515 135
rect 517 133 518 135
rect 514 131 518 133
rect 577 134 587 135
rect 577 132 583 134
rect 585 132 587 134
rect 577 131 587 132
rect 592 134 613 135
rect 592 132 593 134
rect 595 133 613 134
rect 615 133 617 135
rect 622 134 626 136
rect 595 132 617 133
rect 421 118 425 123
rect 452 119 456 130
rect 421 116 422 118
rect 424 116 425 118
rect 421 110 425 116
rect 430 118 456 119
rect 430 116 432 118
rect 434 116 456 118
rect 430 115 456 116
rect 473 119 477 131
rect 504 127 508 131
rect 525 127 529 129
rect 421 109 439 110
rect 421 107 435 109
rect 437 107 439 109
rect 421 106 439 107
rect 433 102 439 106
rect 433 100 435 102
rect 437 100 439 102
rect 433 99 439 100
rect 399 96 403 98
rect 399 94 400 96
rect 402 94 403 96
rect 443 95 447 115
rect 470 118 477 119
rect 470 116 472 118
rect 474 116 477 118
rect 470 115 477 116
rect 473 103 477 115
rect 481 123 508 127
rect 481 118 485 123
rect 481 116 482 118
rect 484 116 485 118
rect 481 111 485 116
rect 490 118 505 119
rect 490 116 492 118
rect 494 116 505 118
rect 490 115 505 116
rect 481 109 498 111
rect 481 107 495 109
rect 497 107 498 109
rect 473 102 489 103
rect 473 100 485 102
rect 487 100 489 102
rect 473 99 489 100
rect 494 102 498 107
rect 494 100 495 102
rect 497 100 498 102
rect 494 98 498 100
rect 501 102 505 115
rect 525 125 526 127
rect 528 125 529 127
rect 525 111 529 125
rect 515 107 529 111
rect 515 102 519 107
rect 501 100 516 102
rect 518 100 519 102
rect 501 98 519 100
rect 577 127 581 131
rect 561 123 581 127
rect 561 120 565 123
rect 559 118 565 120
rect 559 116 560 118
rect 562 116 565 118
rect 559 114 565 116
rect 561 103 565 114
rect 569 118 573 120
rect 592 127 596 132
rect 592 125 593 127
rect 595 125 596 127
rect 592 123 596 125
rect 601 127 616 128
rect 601 125 603 127
rect 605 126 616 127
rect 605 125 630 126
rect 601 124 626 125
rect 612 123 626 124
rect 628 123 630 125
rect 612 122 630 123
rect 569 116 570 118
rect 572 116 573 118
rect 569 111 573 116
rect 612 111 616 122
rect 609 107 616 111
rect 619 115 623 117
rect 619 113 620 115
rect 622 113 623 115
rect 609 106 613 107
rect 609 104 610 106
rect 612 104 613 106
rect 561 102 601 103
rect 609 102 613 104
rect 619 103 623 113
rect 561 100 575 102
rect 577 100 601 102
rect 561 99 601 100
rect 617 99 623 103
rect 501 95 505 98
rect 574 95 578 99
rect 597 95 621 99
rect 370 93 394 94
rect 370 91 390 93
rect 392 91 394 93
rect 370 90 394 91
rect 361 86 363 88
rect 365 86 367 88
rect 361 85 367 86
rect 399 88 403 94
rect 413 94 459 95
rect 413 92 415 94
rect 417 92 455 94
rect 457 92 459 94
rect 413 91 459 92
rect 463 94 469 95
rect 463 92 465 94
rect 467 92 469 94
rect 399 86 400 88
rect 402 86 403 88
rect 399 85 403 86
rect 443 87 449 88
rect 443 85 445 87
rect 447 85 449 87
rect 463 87 469 92
rect 473 94 505 95
rect 473 92 475 94
rect 477 92 505 94
rect 473 91 505 92
rect 524 94 530 95
rect 524 92 526 94
rect 528 92 530 94
rect 463 85 465 87
rect 467 85 469 87
rect 503 87 509 88
rect 503 85 505 87
rect 507 85 509 87
rect 524 85 530 92
rect 563 94 569 95
rect 563 92 565 94
rect 567 92 569 94
rect 563 87 569 92
rect 574 93 575 95
rect 577 93 578 95
rect 574 91 578 93
rect 585 94 591 95
rect 585 92 587 94
rect 589 92 591 94
rect 563 85 565 87
rect 567 85 569 87
rect 585 87 591 92
rect 585 85 587 87
rect 589 85 591 87
rect 620 87 626 88
rect 620 85 622 87
rect 624 85 626 87
rect -182 60 -176 69
rect -182 58 -180 60
rect -178 58 -176 60
rect -182 57 -176 58
rect -171 62 -167 64
rect -171 60 -170 62
rect -168 60 -167 62
rect -171 55 -167 60
rect -162 62 -156 69
rect -162 60 -160 62
rect -158 60 -156 62
rect -162 59 -156 60
rect -137 62 -131 69
rect -111 68 -105 69
rect -111 66 -109 68
rect -107 66 -105 68
rect -137 60 -135 62
rect -133 60 -131 62
rect -137 59 -131 60
rect -120 62 -116 64
rect -120 60 -119 62
rect -117 60 -116 62
rect -171 54 -170 55
rect -184 53 -170 54
rect -168 53 -167 55
rect -184 50 -167 53
rect -184 38 -180 50
rect -120 55 -116 60
rect -111 61 -105 66
rect -73 68 -69 69
rect -73 66 -72 68
rect -70 66 -69 68
rect -29 67 -27 69
rect -25 67 -23 69
rect -29 66 -23 67
rect -9 67 -7 69
rect -5 67 -3 69
rect -111 59 -109 61
rect -107 59 -105 61
rect -111 58 -105 59
rect -102 63 -78 64
rect -102 61 -82 63
rect -80 61 -78 63
rect -102 60 -78 61
rect -73 60 -69 66
rect -102 55 -98 60
rect -73 58 -72 60
rect -70 58 -69 60
rect -59 62 -13 63
rect -59 60 -57 62
rect -55 60 -17 62
rect -15 60 -13 62
rect -59 59 -13 60
rect -9 62 -3 67
rect 31 67 33 69
rect 35 67 37 69
rect 31 66 37 67
rect -9 60 -7 62
rect -5 60 -3 62
rect -9 59 -3 60
rect 1 62 33 63
rect 1 60 3 62
rect 5 60 33 62
rect 1 59 33 60
rect 52 62 58 69
rect 52 60 54 62
rect 56 60 58 62
rect 52 59 58 60
rect 81 62 87 69
rect 107 68 113 69
rect 107 66 109 68
rect 111 66 113 68
rect 81 60 83 62
rect 85 60 87 62
rect 81 59 87 60
rect 98 62 102 64
rect 98 60 99 62
rect 101 60 102 62
rect -73 56 -69 58
rect -120 53 -119 55
rect -117 53 -98 55
rect -120 51 -98 53
rect -184 36 -183 38
rect -181 36 -180 38
rect -184 31 -180 36
rect -184 27 -172 31
rect -188 24 -187 26
rect -176 23 -172 27
rect -144 43 -143 50
rect -39 54 -33 55
rect -39 52 -37 54
rect -35 52 -33 54
rect -176 22 -156 23
rect -176 20 -160 22
rect -158 20 -156 22
rect -176 19 -156 20
rect -144 25 -143 31
rect -133 26 -129 28
rect -133 24 -132 26
rect -130 24 -129 26
rect -133 13 -129 24
rect -85 23 -79 24
rect -85 22 -83 23
rect -124 21 -83 22
rect -81 21 -79 23
rect -124 19 -122 21
rect -120 19 -79 21
rect -124 18 -79 19
rect -75 23 -69 24
rect -75 21 -73 23
rect -71 21 -69 23
rect -75 13 -69 21
rect -39 48 -33 52
rect -51 47 -33 48
rect -51 45 -37 47
rect -35 45 -33 47
rect -51 44 -33 45
rect -51 38 -47 44
rect -29 39 -25 59
rect 29 56 33 59
rect -51 36 -50 38
rect -48 36 -47 38
rect -51 31 -47 36
rect -42 38 -16 39
rect -42 36 -40 38
rect -38 36 -16 38
rect -42 35 -16 36
rect -51 27 -26 31
rect -30 23 -26 27
rect -30 21 -29 23
rect -27 21 -26 23
rect -30 19 -26 21
rect -20 24 -16 35
rect 1 54 17 55
rect 1 52 13 54
rect 15 52 17 54
rect 1 51 17 52
rect 22 54 26 56
rect 22 52 23 54
rect 25 52 26 54
rect 1 39 5 51
rect 22 47 26 52
rect -2 38 5 39
rect -2 36 0 38
rect 2 36 5 38
rect -2 35 5 36
rect -20 23 -3 24
rect -20 21 -7 23
rect -5 21 -3 23
rect -20 20 -3 21
rect 1 23 5 35
rect 9 45 23 47
rect 25 45 26 47
rect 9 43 26 45
rect 29 54 47 56
rect 29 52 44 54
rect 46 52 47 54
rect 9 38 13 43
rect 29 39 33 52
rect 43 47 47 52
rect 43 43 57 47
rect 9 36 10 38
rect 12 36 13 38
rect 9 31 13 36
rect 18 38 33 39
rect 18 36 20 38
rect 22 36 33 38
rect 18 35 33 36
rect 9 27 36 31
rect 53 29 57 43
rect 98 55 102 60
rect 107 61 113 66
rect 145 68 149 69
rect 145 66 146 68
rect 148 66 149 68
rect 189 67 191 69
rect 193 67 195 69
rect 189 66 195 67
rect 209 67 211 69
rect 213 67 215 69
rect 107 59 109 61
rect 111 59 113 61
rect 107 58 113 59
rect 116 63 140 64
rect 116 61 136 63
rect 138 61 140 63
rect 116 60 140 61
rect 145 60 149 66
rect 116 55 120 60
rect 145 58 146 60
rect 148 58 149 60
rect 159 62 205 63
rect 159 60 161 62
rect 163 60 201 62
rect 203 60 205 62
rect 159 59 205 60
rect 209 62 215 67
rect 249 67 251 69
rect 253 67 255 69
rect 249 66 255 67
rect 209 60 211 62
rect 213 60 215 62
rect 209 59 215 60
rect 219 62 251 63
rect 219 60 221 62
rect 223 60 251 62
rect 219 59 251 60
rect 270 62 276 69
rect 270 60 272 62
rect 274 60 276 62
rect 270 59 276 60
rect 301 62 307 69
rect 327 68 333 69
rect 327 66 329 68
rect 331 66 333 68
rect 301 60 303 62
rect 305 60 307 62
rect 301 59 307 60
rect 318 62 322 64
rect 318 60 319 62
rect 321 60 322 62
rect 145 56 149 58
rect 98 53 99 55
rect 101 53 120 55
rect 98 51 120 53
rect 53 27 54 29
rect 56 27 57 29
rect 32 23 36 27
rect 53 25 57 27
rect 74 43 75 50
rect 179 54 185 55
rect 179 52 181 54
rect 183 52 185 54
rect 1 22 27 23
rect 1 20 23 22
rect 25 20 27 22
rect 1 19 27 20
rect 32 21 33 23
rect 35 21 36 23
rect 32 19 36 21
rect 42 21 46 23
rect 42 19 43 21
rect 45 19 46 21
rect -20 15 -14 16
rect -20 13 -18 15
rect -16 13 -14 15
rect 42 13 46 19
rect 74 25 75 31
rect 85 26 89 28
rect 85 24 86 26
rect 88 24 89 26
rect 85 13 89 24
rect 133 23 139 24
rect 133 22 135 23
rect 94 21 135 22
rect 137 21 139 23
rect 94 19 96 21
rect 98 19 139 21
rect 94 18 139 19
rect 143 23 149 24
rect 143 21 145 23
rect 147 21 149 23
rect 143 13 149 21
rect 179 48 185 52
rect 167 47 185 48
rect 167 45 181 47
rect 183 45 185 47
rect 167 44 185 45
rect 167 38 171 44
rect 189 39 193 59
rect 247 56 251 59
rect 167 36 168 38
rect 170 36 171 38
rect 167 31 171 36
rect 176 38 202 39
rect 176 36 178 38
rect 180 36 202 38
rect 176 35 202 36
rect 167 27 192 31
rect 188 23 192 27
rect 188 21 189 23
rect 191 21 192 23
rect 188 19 192 21
rect 198 24 202 35
rect 219 54 235 55
rect 219 52 231 54
rect 233 52 235 54
rect 219 51 235 52
rect 240 54 244 56
rect 240 52 241 54
rect 243 52 244 54
rect 219 39 223 51
rect 240 47 244 52
rect 216 38 223 39
rect 216 36 218 38
rect 220 36 223 38
rect 216 35 223 36
rect 198 23 215 24
rect 198 21 211 23
rect 213 21 215 23
rect 198 20 215 21
rect 219 23 223 35
rect 227 45 241 47
rect 243 45 244 47
rect 227 43 244 45
rect 247 54 265 56
rect 247 52 262 54
rect 264 52 265 54
rect 227 38 231 43
rect 247 39 251 52
rect 261 47 265 52
rect 261 43 275 47
rect 227 36 228 38
rect 230 36 231 38
rect 227 31 231 36
rect 236 38 251 39
rect 236 36 238 38
rect 240 36 251 38
rect 236 35 251 36
rect 227 27 254 31
rect 271 29 275 43
rect 318 55 322 60
rect 327 61 333 66
rect 365 68 369 69
rect 365 66 366 68
rect 368 66 369 68
rect 409 67 411 69
rect 413 67 415 69
rect 409 66 415 67
rect 429 67 431 69
rect 433 67 435 69
rect 327 59 329 61
rect 331 59 333 61
rect 327 58 333 59
rect 336 63 360 64
rect 336 61 356 63
rect 358 61 360 63
rect 336 60 360 61
rect 365 60 369 66
rect 336 55 340 60
rect 365 58 366 60
rect 368 58 369 60
rect 379 62 425 63
rect 379 60 381 62
rect 383 60 421 62
rect 423 60 425 62
rect 379 59 425 60
rect 429 62 435 67
rect 469 67 471 69
rect 473 67 475 69
rect 469 66 475 67
rect 429 60 431 62
rect 433 60 435 62
rect 429 59 435 60
rect 439 62 471 63
rect 439 60 441 62
rect 443 60 471 62
rect 439 59 471 60
rect 490 62 496 69
rect 490 60 492 62
rect 494 60 496 62
rect 490 59 496 60
rect 522 67 524 69
rect 526 67 528 69
rect 522 62 528 67
rect 544 67 546 69
rect 548 67 550 69
rect 522 60 524 62
rect 526 60 528 62
rect 522 59 528 60
rect 533 61 537 63
rect 533 59 534 61
rect 536 59 537 61
rect 544 62 550 67
rect 579 67 581 69
rect 583 67 585 69
rect 579 66 585 67
rect 544 60 546 62
rect 548 60 550 62
rect 544 59 550 60
rect 365 56 369 58
rect 318 53 319 55
rect 321 53 340 55
rect 318 51 340 53
rect 271 27 272 29
rect 274 27 275 29
rect 250 23 254 27
rect 271 25 275 27
rect 294 43 295 50
rect 399 54 405 55
rect 399 52 401 54
rect 403 52 405 54
rect 219 22 245 23
rect 219 20 241 22
rect 243 20 245 22
rect 219 19 245 20
rect 250 21 251 23
rect 253 21 254 23
rect 250 19 254 21
rect 260 21 264 23
rect 260 19 261 21
rect 263 19 264 21
rect 198 15 204 16
rect 198 13 200 15
rect 202 13 204 15
rect 260 13 264 19
rect 294 25 295 31
rect 305 26 309 28
rect 305 24 306 26
rect 308 24 309 26
rect 305 13 309 24
rect 353 23 359 24
rect 353 22 355 23
rect 314 21 355 22
rect 357 21 359 23
rect 314 19 316 21
rect 318 19 359 21
rect 314 18 359 19
rect 363 23 369 24
rect 363 21 365 23
rect 367 21 369 23
rect 363 13 369 21
rect 399 48 405 52
rect 387 47 405 48
rect 387 45 401 47
rect 403 45 405 47
rect 387 44 405 45
rect 387 38 391 44
rect 409 39 413 59
rect 467 56 471 59
rect 387 36 388 38
rect 390 36 391 38
rect 387 31 391 36
rect 396 38 422 39
rect 396 36 398 38
rect 400 36 422 38
rect 396 35 422 36
rect 387 27 412 31
rect 408 23 412 27
rect 408 21 409 23
rect 411 21 412 23
rect 408 19 412 21
rect 418 24 422 35
rect 439 54 455 55
rect 439 52 451 54
rect 453 52 455 54
rect 439 51 455 52
rect 460 54 464 56
rect 460 52 461 54
rect 463 52 464 54
rect 439 39 443 51
rect 460 47 464 52
rect 436 38 443 39
rect 436 36 438 38
rect 440 36 443 38
rect 436 35 443 36
rect 418 23 435 24
rect 418 21 431 23
rect 433 21 435 23
rect 418 20 435 21
rect 439 23 443 35
rect 447 45 461 47
rect 463 45 464 47
rect 447 43 464 45
rect 467 54 485 56
rect 467 52 482 54
rect 484 52 485 54
rect 447 38 451 43
rect 467 39 471 52
rect 481 47 485 52
rect 481 43 495 47
rect 447 36 448 38
rect 450 36 451 38
rect 447 31 451 36
rect 456 38 471 39
rect 456 36 458 38
rect 460 36 471 38
rect 456 35 471 36
rect 447 27 474 31
rect 491 29 495 43
rect 533 55 537 59
rect 556 55 580 59
rect 520 54 560 55
rect 520 52 534 54
rect 536 52 560 54
rect 520 51 560 52
rect 491 27 492 29
rect 494 27 495 29
rect 470 23 474 27
rect 491 25 495 27
rect 520 40 524 51
rect 568 50 572 52
rect 576 51 582 55
rect 568 48 569 50
rect 571 48 572 50
rect 568 47 572 48
rect 568 43 575 47
rect 518 38 524 40
rect 518 36 519 38
rect 521 36 524 38
rect 518 34 524 36
rect 528 38 532 43
rect 528 36 529 38
rect 531 36 532 38
rect 528 34 532 36
rect 520 31 524 34
rect 520 27 540 31
rect 536 23 540 27
rect 571 32 575 43
rect 578 41 582 51
rect 578 39 579 41
rect 581 39 582 41
rect 578 37 582 39
rect 571 31 589 32
rect 551 29 555 31
rect 571 30 585 31
rect 551 27 552 29
rect 554 27 555 29
rect 439 22 465 23
rect 439 20 461 22
rect 463 20 465 22
rect 439 19 465 20
rect 470 21 471 23
rect 473 21 474 23
rect 470 19 474 21
rect 480 21 484 23
rect 480 19 481 21
rect 483 19 484 21
rect 536 22 546 23
rect 536 20 542 22
rect 544 20 546 22
rect 536 19 546 20
rect 551 22 555 27
rect 560 29 585 30
rect 587 29 589 31
rect 560 27 562 29
rect 564 28 589 29
rect 564 27 575 28
rect 560 26 575 27
rect 551 20 552 22
rect 554 21 576 22
rect 554 20 572 21
rect 551 19 572 20
rect 574 19 576 21
rect 418 15 424 16
rect 418 13 420 15
rect 422 13 424 15
rect 480 13 484 19
rect 551 18 576 19
rect 581 18 585 20
rect 581 16 582 18
rect 584 16 585 18
rect 523 15 529 16
rect 523 13 525 15
rect 527 13 529 15
rect 581 13 585 16
rect -195 -14 -191 -3
rect -186 -9 -141 -8
rect -186 -11 -184 -9
rect -182 -11 -141 -9
rect -186 -12 -145 -11
rect -147 -13 -145 -12
rect -143 -13 -141 -11
rect -147 -14 -141 -13
rect -137 -11 -131 -3
rect -82 -5 -80 -3
rect -78 -5 -76 -3
rect -82 -6 -76 -5
rect -20 -9 -16 -3
rect -137 -13 -135 -11
rect -133 -13 -131 -11
rect -137 -14 -131 -13
rect -92 -11 -88 -9
rect -61 -10 -35 -9
rect -92 -13 -91 -11
rect -89 -13 -88 -11
rect -206 -21 -205 -15
rect -195 -16 -194 -14
rect -192 -16 -191 -14
rect -195 -18 -191 -16
rect -206 -40 -205 -33
rect -182 -43 -160 -41
rect -182 -45 -181 -43
rect -179 -45 -160 -43
rect -199 -50 -193 -49
rect -199 -52 -197 -50
rect -195 -52 -193 -50
rect -199 -59 -193 -52
rect -182 -50 -178 -45
rect -182 -52 -181 -50
rect -179 -52 -178 -50
rect -182 -54 -178 -52
rect -173 -49 -167 -48
rect -173 -51 -171 -49
rect -169 -51 -167 -49
rect -173 -56 -167 -51
rect -164 -50 -160 -45
rect -92 -17 -88 -13
rect -113 -21 -88 -17
rect -82 -11 -65 -10
rect -82 -13 -69 -11
rect -67 -13 -65 -11
rect -82 -14 -65 -13
rect -61 -12 -39 -10
rect -37 -12 -35 -10
rect -61 -13 -35 -12
rect -30 -11 -26 -9
rect -30 -13 -29 -11
rect -27 -13 -26 -11
rect -20 -11 -19 -9
rect -17 -11 -16 -9
rect -20 -13 -16 -11
rect -113 -26 -109 -21
rect -82 -25 -78 -14
rect -113 -28 -112 -26
rect -110 -28 -109 -26
rect -113 -34 -109 -28
rect -104 -26 -78 -25
rect -104 -28 -102 -26
rect -100 -28 -78 -26
rect -104 -29 -78 -28
rect -61 -25 -57 -13
rect -30 -17 -26 -13
rect -9 -17 -5 -15
rect -113 -35 -95 -34
rect -113 -37 -99 -35
rect -97 -37 -95 -35
rect -113 -38 -95 -37
rect -101 -42 -95 -38
rect -101 -44 -99 -42
rect -97 -44 -95 -42
rect -101 -45 -95 -44
rect -135 -48 -131 -46
rect -135 -50 -134 -48
rect -132 -50 -131 -48
rect -91 -49 -87 -29
rect -64 -26 -57 -25
rect -64 -28 -62 -26
rect -60 -28 -57 -26
rect -64 -29 -57 -28
rect -61 -41 -57 -29
rect -53 -21 -26 -17
rect -53 -26 -49 -21
rect -53 -28 -52 -26
rect -50 -28 -49 -26
rect -53 -33 -49 -28
rect -44 -26 -29 -25
rect -44 -28 -42 -26
rect -40 -28 -29 -26
rect -44 -29 -29 -28
rect -53 -35 -36 -33
rect -53 -37 -39 -35
rect -37 -37 -36 -35
rect -61 -42 -45 -41
rect -61 -44 -49 -42
rect -47 -44 -45 -42
rect -61 -45 -45 -44
rect -40 -42 -36 -37
rect -40 -44 -39 -42
rect -37 -44 -36 -42
rect -40 -46 -36 -44
rect -33 -42 -29 -29
rect -9 -19 -8 -17
rect -6 -19 -5 -17
rect -9 -33 -5 -19
rect 25 -14 29 -3
rect 34 -9 79 -8
rect 34 -11 36 -9
rect 38 -11 79 -9
rect 34 -12 75 -11
rect 73 -13 75 -12
rect 77 -13 79 -11
rect 73 -14 79 -13
rect 83 -11 89 -3
rect 138 -5 140 -3
rect 142 -5 144 -3
rect 138 -6 144 -5
rect 200 -9 204 -3
rect 83 -13 85 -11
rect 87 -13 89 -11
rect 83 -14 89 -13
rect 128 -11 132 -9
rect 159 -10 185 -9
rect 128 -13 129 -11
rect 131 -13 132 -11
rect -19 -37 -5 -33
rect -19 -42 -15 -37
rect -33 -44 -18 -42
rect -16 -44 -15 -42
rect -33 -46 -15 -44
rect 14 -21 15 -15
rect 25 -16 26 -14
rect 28 -16 29 -14
rect 25 -18 29 -16
rect 14 -40 15 -33
rect 38 -43 60 -41
rect 38 -45 39 -43
rect 41 -45 60 -43
rect -33 -49 -29 -46
rect -164 -51 -140 -50
rect -164 -53 -144 -51
rect -142 -53 -140 -51
rect -164 -54 -140 -53
rect -173 -58 -171 -56
rect -169 -58 -167 -56
rect -173 -59 -167 -58
rect -135 -56 -131 -50
rect -121 -50 -75 -49
rect -121 -52 -119 -50
rect -117 -52 -79 -50
rect -77 -52 -75 -50
rect -121 -53 -75 -52
rect -71 -50 -65 -49
rect -71 -52 -69 -50
rect -67 -52 -65 -50
rect -135 -58 -134 -56
rect -132 -58 -131 -56
rect -135 -59 -131 -58
rect -91 -57 -85 -56
rect -91 -59 -89 -57
rect -87 -59 -85 -57
rect -71 -57 -65 -52
rect -61 -50 -29 -49
rect -61 -52 -59 -50
rect -57 -52 -29 -50
rect -61 -53 -29 -52
rect -10 -50 -4 -49
rect -10 -52 -8 -50
rect -6 -52 -4 -50
rect -71 -59 -69 -57
rect -67 -59 -65 -57
rect -31 -57 -25 -56
rect -31 -59 -29 -57
rect -27 -59 -25 -57
rect -10 -59 -4 -52
rect 21 -50 27 -49
rect 21 -52 23 -50
rect 25 -52 27 -50
rect 21 -59 27 -52
rect 38 -50 42 -45
rect 38 -52 39 -50
rect 41 -52 42 -50
rect 38 -54 42 -52
rect 47 -49 53 -48
rect 47 -51 49 -49
rect 51 -51 53 -49
rect 47 -56 53 -51
rect 56 -50 60 -45
rect 128 -17 132 -13
rect 107 -21 132 -17
rect 138 -11 155 -10
rect 138 -13 151 -11
rect 153 -13 155 -11
rect 138 -14 155 -13
rect 159 -12 181 -10
rect 183 -12 185 -10
rect 159 -13 185 -12
rect 190 -11 194 -9
rect 190 -13 191 -11
rect 193 -13 194 -11
rect 200 -11 201 -9
rect 203 -11 204 -9
rect 200 -13 204 -11
rect 107 -26 111 -21
rect 138 -25 142 -14
rect 107 -28 108 -26
rect 110 -28 111 -26
rect 107 -34 111 -28
rect 116 -26 142 -25
rect 116 -28 118 -26
rect 120 -28 142 -26
rect 116 -29 142 -28
rect 159 -25 163 -13
rect 190 -17 194 -13
rect 211 -17 215 -15
rect 107 -35 125 -34
rect 107 -37 121 -35
rect 123 -37 125 -35
rect 107 -38 125 -37
rect 119 -42 125 -38
rect 119 -44 121 -42
rect 123 -44 125 -42
rect 119 -45 125 -44
rect 85 -48 89 -46
rect 85 -50 86 -48
rect 88 -50 89 -48
rect 129 -49 133 -29
rect 156 -26 163 -25
rect 156 -28 158 -26
rect 160 -28 163 -26
rect 156 -29 163 -28
rect 159 -41 163 -29
rect 167 -21 194 -17
rect 167 -26 171 -21
rect 167 -28 168 -26
rect 170 -28 171 -26
rect 167 -33 171 -28
rect 176 -26 191 -25
rect 176 -28 178 -26
rect 180 -28 191 -26
rect 176 -29 191 -28
rect 167 -35 184 -33
rect 167 -37 181 -35
rect 183 -37 184 -35
rect 159 -42 175 -41
rect 159 -44 171 -42
rect 173 -44 175 -42
rect 159 -45 175 -44
rect 180 -42 184 -37
rect 180 -44 181 -42
rect 183 -44 184 -42
rect 180 -46 184 -44
rect 187 -42 191 -29
rect 211 -19 212 -17
rect 214 -19 215 -17
rect 211 -33 215 -19
rect 242 -14 246 -3
rect 251 -9 296 -8
rect 251 -11 253 -9
rect 255 -11 296 -9
rect 251 -12 292 -11
rect 290 -13 292 -12
rect 294 -13 296 -11
rect 290 -14 296 -13
rect 300 -11 306 -3
rect 355 -5 357 -3
rect 359 -5 361 -3
rect 355 -6 361 -5
rect 417 -9 421 -3
rect 466 -5 468 -3
rect 470 -5 472 -3
rect 466 -6 472 -5
rect 524 -6 528 -3
rect 524 -8 525 -6
rect 527 -8 528 -6
rect 494 -9 519 -8
rect 300 -13 302 -11
rect 304 -13 306 -11
rect 300 -14 306 -13
rect 345 -11 349 -9
rect 376 -10 402 -9
rect 345 -13 346 -11
rect 348 -13 349 -11
rect 201 -37 215 -33
rect 201 -42 205 -37
rect 187 -44 202 -42
rect 204 -44 205 -42
rect 187 -46 205 -44
rect 231 -21 232 -15
rect 242 -16 243 -14
rect 245 -16 246 -14
rect 242 -18 246 -16
rect 231 -40 232 -33
rect 255 -43 277 -41
rect 255 -45 256 -43
rect 258 -45 277 -43
rect 187 -49 191 -46
rect 56 -51 80 -50
rect 56 -53 76 -51
rect 78 -53 80 -51
rect 56 -54 80 -53
rect 47 -58 49 -56
rect 51 -58 53 -56
rect 47 -59 53 -58
rect 85 -56 89 -50
rect 99 -50 145 -49
rect 99 -52 101 -50
rect 103 -52 141 -50
rect 143 -52 145 -50
rect 99 -53 145 -52
rect 149 -50 155 -49
rect 149 -52 151 -50
rect 153 -52 155 -50
rect 85 -58 86 -56
rect 88 -58 89 -56
rect 85 -59 89 -58
rect 129 -57 135 -56
rect 129 -59 131 -57
rect 133 -59 135 -57
rect 149 -57 155 -52
rect 159 -50 191 -49
rect 159 -52 161 -50
rect 163 -52 191 -50
rect 159 -53 191 -52
rect 210 -50 216 -49
rect 210 -52 212 -50
rect 214 -52 216 -50
rect 149 -59 151 -57
rect 153 -59 155 -57
rect 189 -57 195 -56
rect 189 -59 191 -57
rect 193 -59 195 -57
rect 210 -59 216 -52
rect 238 -50 244 -49
rect 238 -52 240 -50
rect 242 -52 244 -50
rect 238 -59 244 -52
rect 255 -50 259 -45
rect 255 -52 256 -50
rect 258 -52 259 -50
rect 255 -54 259 -52
rect 264 -49 270 -48
rect 264 -51 266 -49
rect 268 -51 270 -49
rect 264 -56 270 -51
rect 273 -50 277 -45
rect 345 -17 349 -13
rect 324 -21 349 -17
rect 355 -11 372 -10
rect 355 -13 368 -11
rect 370 -13 372 -11
rect 355 -14 372 -13
rect 376 -12 398 -10
rect 400 -12 402 -10
rect 376 -13 402 -12
rect 407 -11 411 -9
rect 407 -13 408 -11
rect 410 -13 411 -11
rect 417 -11 418 -9
rect 420 -11 421 -9
rect 417 -13 421 -11
rect 479 -10 489 -9
rect 479 -12 485 -10
rect 487 -12 489 -10
rect 479 -13 489 -12
rect 494 -10 515 -9
rect 494 -12 495 -10
rect 497 -11 515 -10
rect 517 -11 519 -9
rect 524 -10 528 -8
rect 497 -12 519 -11
rect 324 -26 328 -21
rect 355 -25 359 -14
rect 324 -28 325 -26
rect 327 -28 328 -26
rect 324 -34 328 -28
rect 333 -26 359 -25
rect 333 -28 335 -26
rect 337 -28 359 -26
rect 333 -29 359 -28
rect 376 -25 380 -13
rect 407 -17 411 -13
rect 428 -17 432 -15
rect 324 -35 342 -34
rect 324 -37 338 -35
rect 340 -37 342 -35
rect 324 -38 342 -37
rect 336 -42 342 -38
rect 336 -44 338 -42
rect 340 -44 342 -42
rect 336 -45 342 -44
rect 302 -48 306 -46
rect 302 -50 303 -48
rect 305 -50 306 -48
rect 346 -49 350 -29
rect 373 -26 380 -25
rect 373 -28 375 -26
rect 377 -28 380 -26
rect 373 -29 380 -28
rect 376 -41 380 -29
rect 384 -21 411 -17
rect 384 -26 388 -21
rect 384 -28 385 -26
rect 387 -28 388 -26
rect 384 -33 388 -28
rect 393 -26 408 -25
rect 393 -28 395 -26
rect 397 -28 408 -26
rect 393 -29 408 -28
rect 384 -35 401 -33
rect 384 -37 398 -35
rect 400 -37 401 -35
rect 376 -42 392 -41
rect 376 -44 388 -42
rect 390 -44 392 -42
rect 376 -45 392 -44
rect 397 -42 401 -37
rect 397 -44 398 -42
rect 400 -44 401 -42
rect 397 -46 401 -44
rect 404 -42 408 -29
rect 428 -19 429 -17
rect 431 -19 432 -17
rect 428 -33 432 -19
rect 418 -37 432 -33
rect 418 -42 422 -37
rect 404 -44 419 -42
rect 421 -44 422 -42
rect 404 -46 422 -44
rect 479 -17 483 -13
rect 463 -21 483 -17
rect 463 -24 467 -21
rect 461 -26 467 -24
rect 461 -28 462 -26
rect 464 -28 467 -26
rect 461 -30 467 -28
rect 463 -41 467 -30
rect 471 -26 475 -24
rect 494 -17 498 -12
rect 494 -19 495 -17
rect 497 -19 498 -17
rect 494 -21 498 -19
rect 503 -17 518 -16
rect 503 -19 505 -17
rect 507 -18 518 -17
rect 507 -19 532 -18
rect 503 -20 528 -19
rect 514 -21 528 -20
rect 530 -21 532 -19
rect 514 -22 532 -21
rect 471 -28 472 -26
rect 474 -28 475 -26
rect 471 -33 475 -28
rect 514 -33 518 -22
rect 511 -37 518 -33
rect 521 -29 525 -27
rect 521 -31 522 -29
rect 524 -31 525 -29
rect 511 -38 515 -37
rect 511 -40 512 -38
rect 514 -40 515 -38
rect 463 -42 503 -41
rect 511 -42 515 -40
rect 521 -41 525 -31
rect 463 -44 477 -42
rect 479 -44 503 -42
rect 463 -45 503 -44
rect 519 -45 525 -41
rect 404 -49 408 -46
rect 476 -49 480 -45
rect 499 -49 523 -45
rect 273 -51 297 -50
rect 273 -53 293 -51
rect 295 -53 297 -51
rect 273 -54 297 -53
rect 264 -58 266 -56
rect 268 -58 270 -56
rect 264 -59 270 -58
rect 302 -56 306 -50
rect 316 -50 362 -49
rect 316 -52 318 -50
rect 320 -52 358 -50
rect 360 -52 362 -50
rect 316 -53 362 -52
rect 366 -50 372 -49
rect 366 -52 368 -50
rect 370 -52 372 -50
rect 302 -58 303 -56
rect 305 -58 306 -56
rect 302 -59 306 -58
rect 346 -57 352 -56
rect 346 -59 348 -57
rect 350 -59 352 -57
rect 366 -57 372 -52
rect 376 -50 408 -49
rect 376 -52 378 -50
rect 380 -52 408 -50
rect 376 -53 408 -52
rect 427 -50 433 -49
rect 427 -52 429 -50
rect 431 -52 433 -50
rect 366 -59 368 -57
rect 370 -59 372 -57
rect 406 -57 412 -56
rect 406 -59 408 -57
rect 410 -59 412 -57
rect 427 -59 433 -52
rect 465 -50 471 -49
rect 465 -52 467 -50
rect 469 -52 471 -50
rect 465 -57 471 -52
rect 476 -51 477 -49
rect 479 -51 480 -49
rect 476 -53 480 -51
rect 487 -50 493 -49
rect 487 -52 489 -50
rect 491 -52 493 -50
rect 465 -59 467 -57
rect 469 -59 471 -57
rect 487 -57 493 -52
rect 487 -59 489 -57
rect 491 -59 493 -57
rect 522 -57 528 -56
rect 522 -59 524 -57
rect 526 -59 528 -57
<< via1 >>
rect 75 196 77 198
rect 115 196 117 198
rect 67 178 69 180
rect 48 162 50 164
rect 107 179 109 181
rect 84 162 86 164
rect 158 191 160 193
rect 127 162 129 164
rect 151 170 153 172
rect 262 191 264 193
rect 304 196 306 198
rect 234 162 236 164
rect 254 171 256 173
rect 348 196 350 198
rect 296 179 298 181
rect 272 162 274 164
rect 316 171 318 173
rect 417 196 419 198
rect 340 171 342 173
rect 461 196 463 198
rect 388 162 390 164
rect 409 171 411 173
rect 437 163 439 165
rect 453 171 455 173
rect 503 191 505 193
rect 544 195 546 197
rect 495 179 497 181
rect 471 162 473 164
rect 587 196 589 198
rect 519 162 521 164
rect 536 171 538 173
rect 579 179 581 181
rect 562 162 564 164
rect 627 191 629 193
rect 670 196 672 198
rect 602 162 604 164
rect 620 170 622 172
rect 663 170 665 172
rect -74 103 -72 105
rect -59 116 -57 118
rect -42 108 -40 110
rect -32 102 -30 104
rect -17 116 -15 118
rect 48 124 50 126
rect 0 108 2 110
rect 16 103 18 105
rect 64 117 66 119
rect 115 125 117 127
rect 147 124 149 126
rect 180 124 182 126
rect 139 116 141 118
rect 115 100 117 102
rect 87 92 89 94
rect 171 99 173 101
rect 244 119 246 121
rect 200 100 202 102
rect 292 117 294 119
rect 316 117 318 119
rect 308 100 310 102
rect 333 125 335 127
rect 365 124 367 126
rect 388 124 390 126
rect 398 124 400 126
rect 357 116 359 118
rect 333 100 335 102
rect 389 99 391 101
rect 462 119 464 121
rect 421 100 423 102
rect 510 117 512 119
rect 534 117 536 119
rect 526 100 528 102
rect 586 124 588 126
rect 554 104 556 106
rect 602 117 604 119
rect -159 53 -157 55
rect -176 36 -174 38
rect -191 19 -189 21
rect -83 53 -81 55
rect -115 36 -113 38
rect -139 27 -137 29
rect -107 28 -105 30
rect -74 28 -72 30
rect -147 19 -145 21
rect -47 20 -45 22
rect -10 33 -8 35
rect 54 52 56 54
rect 38 35 40 37
rect 135 53 137 55
rect 103 36 105 38
rect 79 27 81 29
rect 111 28 113 30
rect 144 28 146 30
rect 71 19 73 21
rect 170 20 172 22
rect 208 33 210 35
rect 272 52 274 54
rect 256 35 258 37
rect 355 53 357 55
rect 323 36 325 38
rect 299 27 301 29
rect 346 36 348 38
rect 331 28 333 30
rect 364 28 366 30
rect 291 19 293 21
rect 391 20 393 22
rect 428 33 430 35
rect 492 52 494 54
rect 476 35 478 37
rect 553 44 555 46
rect 536 36 538 38
rect 512 23 514 25
rect -201 -19 -199 -17
rect -169 -20 -167 -18
rect -136 -20 -134 -18
rect -177 -28 -175 -26
rect -145 -45 -143 -43
rect -72 -25 -70 -23
rect -24 -27 -22 -25
rect -8 -44 -6 -42
rect 19 -19 21 -17
rect 51 -20 53 -18
rect 84 -20 86 -18
rect 43 -28 45 -26
rect 11 -41 13 -39
rect 75 -45 77 -43
rect 148 -25 150 -23
rect 196 -27 198 -25
rect 212 -44 214 -42
rect 236 -19 238 -17
rect 268 -20 270 -18
rect 291 -20 293 -18
rect 301 -20 303 -18
rect 260 -28 262 -26
rect 228 -40 230 -38
rect 292 -45 294 -43
rect 365 -25 367 -23
rect 413 -27 415 -25
rect 429 -44 431 -42
rect 488 -19 490 -17
rect 455 -41 457 -39
rect 472 -36 474 -34
<< via2 >>
rect -159 211 -157 213
rect -176 148 -174 150
rect -42 211 -40 213
rect -59 159 -57 161
rect 115 211 117 213
rect 0 200 2 202
rect -17 148 -15 150
rect 75 200 77 202
rect 348 211 350 213
rect 304 200 306 202
rect 417 200 419 202
rect 461 200 463 202
rect 544 201 546 203
rect 587 201 589 203
rect 670 201 672 203
rect 158 187 160 189
rect 262 187 264 189
rect 503 187 505 189
rect 627 187 629 189
rect 108 175 110 177
rect 297 175 299 177
rect 67 159 69 161
rect 65 131 67 133
rect 84 131 86 133
rect 115 130 117 132
rect -83 59 -81 61
rect -74 59 -72 61
rect -115 44 -113 46
rect -32 44 -30 46
rect -139 22 -137 24
rect -201 -14 -199 -12
rect -107 22 -105 24
rect -74 24 -72 26
rect -10 26 -8 28
rect 54 59 56 61
rect 39 44 41 46
rect 495 175 497 177
rect 579 175 581 177
rect 150 148 152 150
rect 147 130 149 132
rect 180 128 182 130
rect 255 159 257 161
rect 234 128 236 130
rect 244 126 246 128
rect 139 108 141 110
rect 272 108 274 110
rect 340 167 342 169
rect 409 167 411 169
rect 333 130 335 132
rect 365 130 367 132
rect 398 128 400 130
rect 293 108 295 110
rect 357 108 359 110
rect 171 93 173 95
rect 127 82 129 84
rect 144 82 146 84
rect 115 59 117 61
rect 135 59 137 61
rect 87 44 89 46
rect 103 44 105 46
rect 15 26 17 28
rect 79 22 81 24
rect -169 -14 -167 -12
rect 111 22 113 24
rect 308 93 310 95
rect 200 80 202 82
rect 323 80 325 82
rect 272 59 274 61
rect 257 44 259 46
rect 144 24 146 26
rect 389 93 391 95
rect 421 82 423 84
rect 333 59 335 61
rect 346 59 348 61
rect 323 44 325 46
rect 355 59 357 61
rect 453 149 455 151
rect 462 126 464 128
rect 620 167 622 169
rect 537 159 539 161
rect 663 167 665 169
rect 519 132 521 134
rect 534 132 536 134
rect 471 108 473 110
rect 562 132 564 134
rect 586 132 588 134
rect 511 108 513 110
rect 526 93 528 95
rect 536 82 538 84
rect 437 59 439 61
rect 492 59 494 61
rect 477 44 479 46
rect 208 26 210 28
rect 299 22 301 24
rect -47 7 -45 9
rect 43 7 45 9
rect -147 -16 -145 -14
rect 19 -14 21 -12
rect -136 -16 -134 -14
rect -72 -18 -70 -16
rect -191 -36 -189 -34
rect -177 -36 -175 -34
rect -23 -36 -21 -34
rect 51 -14 53 -12
rect 331 22 333 24
rect 364 24 366 26
rect 428 26 430 28
rect 170 7 172 9
rect 259 7 261 9
rect 71 -16 73 -14
rect 236 -14 238 -12
rect 84 -16 86 -14
rect 148 -18 150 -16
rect 43 -36 45 -34
rect 197 -36 199 -34
rect 268 -14 270 -12
rect 391 7 393 9
rect 471 7 473 9
rect 301 -16 303 -14
rect 365 -18 367 -16
rect 260 -36 262 -34
rect 414 -36 416 -34
rect 488 7 490 9
rect 512 7 514 9
rect -145 -51 -143 -49
rect -8 -51 -6 -49
rect 11 -51 13 -49
rect 75 -51 77 -49
rect 212 -51 214 -49
rect 228 -51 230 -49
rect 292 -51 294 -49
rect 429 -51 431 -49
rect 455 -51 457 -49
<< labels >>
rlabel alu1 612 152 612 152 6 vss
rlabel alu1 612 216 612 216 6 vdd
rlabel alu1 612 180 612 180 1 a0
rlabel alu1 620 176 620 176 1 a0
rlabel alu1 620 188 620 188 1 b1
rlabel alu1 628 196 628 196 1 b1
rlabel alu1 596 180 596 180 1 a0b1
rlabel alu1 604 164 604 164 1 a0b1
rlabel alu1 572 152 572 152 6 vss
rlabel alu1 572 216 572 216 6 vdd
rlabel alu1 572 180 572 180 1 a1
rlabel alu1 580 176 580 176 1 a1
rlabel alu1 580 188 580 188 1 b0
rlabel alu1 556 180 556 180 1 a1b0
rlabel alu1 564 164 564 164 1 a1b0
rlabel alu1 591 81 591 81 2 vdd
rlabel alu1 591 145 591 145 2 vss
rlabel ndifct1 555 133 555 133 1 c01
rlabel alu1 563 133 563 133 1 c01
rlabel alu1 571 133 571 133 1 c01
rlabel via1 555 105 555 105 1 c01
rlabel alu0 582 133 582 133 1 c01_inv
rlabel alu0 563 113 563 113 1 c01_inv
rlabel alu0 576 97 576 97 1 c01_inv
rlabel alu0 581 101 581 101 1 c01_inv
rlabel alu1 635 117 635 117 1 res1
rlabel alu1 627 93 627 93 1 res1
rlabel alu0 621 108 621 108 1 c01_inv
rlabel alu0 621 124 621 124 1 res1_inv
rlabel alu0 611 107 611 107 1 res1_inv
rlabel alu0 609 126 609 126 1 res1_inv
rlabel alu1 587 121 587 121 1 a1b0
rlabel alu1 579 117 579 117 1 a1b0
rlabel alu1 571 109 571 109 1 a0b1
rlabel alu1 579 109 579 109 1 a0b1
rlabel alu1 587 109 587 109 1 a0b1
rlabel alu1 595 109 595 109 1 a0b1
rlabel alu1 603 113 603 113 1 a0b1
rlabel alu1 655 152 655 152 6 vss
rlabel alu1 655 216 655 216 6 vdd
rlabel alu1 655 180 655 180 1 a0
rlabel alu1 663 176 663 176 1 a0
rlabel alu1 663 188 663 188 1 b0
rlabel alu1 588 196 588 196 1 b0
rlabel alu1 671 196 671 196 1 b0
rlabel alu1 639 180 639 180 1 res0
rlabel alu1 647 164 647 164 1 res0
rlabel alu0 663 164 663 164 1 res0_inv
rlabel alu0 647 183 647 183 1 res0_inv
rlabel alu1 475 81 475 81 8 vdd
rlabel alu1 475 145 475 145 8 vss
rlabel alu1 378 81 378 81 8 vdd
rlabel alu1 378 145 378 145 8 vss
rlabel alu1 334 81 334 81 8 vdd
rlabel alu1 334 145 334 145 8 vss
rlabel alu1 326 117 326 117 1 c02
rlabel via1 334 101 334 101 1 c02
rlabel alu1 334 121 334 121 1 c02_inv
rlabel alu1 374 125 374 125 1 c02_inv
rlabel alu1 342 117 342 117 1 c02_inv
rlabel alu1 423 101 423 101 1 s02
rlabel alu1 415 117 415 117 1 s02
rlabel alu1 423 133 423 133 1 s02
rlabel alu1 431 133 431 133 1 s02
rlabel alu0 370 134 370 134 1 fa_11_n3
rlabel alu0 390 133 390 133 1 fa_11_n3
rlabel alu0 354 97 354 97 1 fa_11_n1
rlabel alu0 382 92 382 92 1 fa_11_n1
rlabel alu1 529 152 529 152 6 vss
rlabel alu1 529 216 529 216 6 vdd
rlabel alu1 529 180 529 180 1 a2
rlabel alu1 537 176 537 176 1 a2
rlabel alu1 537 188 537 188 1 b0
rlabel via1 545 196 545 196 1 b0
rlabel alu1 513 180 513 180 1 a2b0
rlabel alu1 521 164 521 164 1 a2b0
rlabel polyct1 535 109 535 109 1 a2b0
rlabel alu1 398 113 398 113 1 a2b0
rlabel alu1 488 216 488 216 6 vdd
rlabel alu1 488 152 488 152 6 vss
rlabel alu1 488 180 488 180 1 a1
rlabel alu1 496 176 496 176 1 a1
rlabel alu1 496 188 496 188 1 b1
rlabel alu1 504 196 504 196 1 b1
rlabel alu1 472 180 472 180 1 a1b1
rlabel alu1 350 113 350 113 1 a1b1
rlabel alu1 519 121 519 121 1 a1b1
rlabel alu1 480 164 480 164 1 a1b1
rlabel alu1 446 152 446 152 6 vss
rlabel alu1 446 216 446 216 6 vdd
rlabel alu1 446 180 446 180 1 a3
rlabel alu1 454 176 454 176 1 a3
rlabel alu1 462 196 462 196 1 b0
rlabel alu1 430 180 430 180 1 a3b0
rlabel via1 438 164 438 164 1 a3b0
rlabel alu0 438 183 438 183 1 a3b0_inv
rlabel alu0 451 200 451 200 1 a3b0_inv
rlabel alu1 454 188 454 188 1 b0
rlabel alu1 402 216 402 216 6 vdd
rlabel alu1 402 152 402 152 6 vss
rlabel alu1 410 188 410 188 1 b2
rlabel alu1 402 180 402 180 1 a0
rlabel alu1 410 176 410 176 1 a0
rlabel alu1 386 180 386 180 1 a0b2
rlabel alu1 394 164 394 164 1 a0b2
rlabel alu1 390 125 390 125 1 a0b2
rlabel alu1 382 117 382 117 1 a0b2
rlabel alu1 463 113 463 113 1 a0b2
rlabel alu1 455 101 455 101 1 a0b2
rlabel alu0 407 200 407 200 1 a0b2_inv_0
rlabel alu0 410 164 410 164 1 a0b2_inv_0
rlabel alu0 496 164 496 164 1 a1b1_inv_0
rlabel alu0 521 183 521 183 1 a2b0_inv_0
rlabel alu0 537 164 537 164 1 a2b0_inv_0
rlabel alu0 564 183 564 183 1 a1b0_inv_0
rlabel alu0 580 164 580 164 1 a1b0_inv_0
rlabel alu0 604 183 604 183 1 a0b1_inv_0
rlabel alu0 620 164 620 164 1 a0b1_inv_0
rlabel alu0 496 105 496 105 1 a1b1_inv_1
rlabel alu0 527 118 527 118 1 a2b0_inv_1
rlabel alu0 517 105 517 105 1 a2b0_inv_1
rlabel alu0 497 117 497 117 1 a2b0_inv_1
rlabel alu0 445 105 445 105 1 a0b2_inv_1
rlabel alu0 480 183 480 183 1 a1b1_inv_0
rlabel alu1 116 145 116 145 8 vss
rlabel alu1 116 81 116 81 8 vdd
rlabel alu1 160 145 160 145 8 vss
rlabel alu1 160 81 160 81 8 vdd
rlabel alu1 257 145 257 145 8 vss
rlabel alu1 257 81 257 81 8 vdd
rlabel alu1 108 117 108 117 1 c03
rlabel via1 116 101 116 101 1 c03
rlabel alu1 116 121 116 121 1 c03_inv
rlabel alu1 124 117 124 117 1 c03_inv
rlabel alu1 156 125 156 125 1 c03_inv
rlabel alu1 213 133 213 133 1 s03
rlabel alu1 205 133 205 133 1 s03
rlabel alu1 197 117 197 117 1 s03
rlabel alu1 205 101 205 101 1 s03
rlabel alu0 152 134 152 134 1 fa_12_n3
rlabel alu0 172 133 172 133 1 fa_12_n3
rlabel alu0 164 92 164 92 1 fa_12_n1
rlabel alu0 136 97 136 97 1 fa_12_n1
rlabel alu1 333 216 333 216 6 vdd
rlabel alu1 333 152 333 152 6 vss
rlabel alu1 349 196 349 196 1 b3
rlabel alu1 341 188 341 188 1 b3
rlabel alu1 333 180 333 180 1 a0
rlabel alu1 341 176 341 176 1 a0
rlabel alu1 317 180 317 180 1 a0b3
rlabel alu1 325 164 325 164 1 a0b3
rlabel alu0 338 200 338 200 1 a0b3_inv_0
rlabel alu0 325 183 325 183 1 a0b3_inv_0
rlabel alu0 341 164 341 164 1 a0b3_inv_0
rlabel polyct1 317 109 317 109 1 a0b3
rlabel alu1 172 104 172 104 1 a0b3
rlabel alu1 180 113 180 113 1 a0b3
rlabel alu0 309 118 309 118 1 a0b3_inv_1
rlabel alu0 299 105 299 105 1 a0b3_inv_1
rlabel alu0 279 117 279 117 1 a0b3_inv_1
rlabel alu1 289 216 289 216 6 vdd
rlabel alu1 289 152 289 152 6 vss
rlabel alu1 305 196 305 196 1 b2
rlabel alu1 297 188 297 188 1 b2
rlabel alu1 289 180 289 180 1 a1
rlabel alu1 297 176 297 176 1 a1
rlabel alu1 418 196 418 196 1 b2
rlabel alu1 273 180 273 180 1 a1b2
rlabel alu1 281 164 281 164 1 a1b2
rlabel alu0 294 200 294 200 1 a1b2_inv_0
rlabel alu0 281 183 281 183 1 a1b2_inv_0
rlabel alu0 297 164 297 164 1 a1b2_inv_0
rlabel alu1 301 121 301 121 1 a1b2
rlabel alu1 132 113 132 113 1 a1b2
rlabel alu0 288 129 288 129 1 a1b2_inv_1
rlabel polyct0 265 117 265 117 1 a1b2_inv_1
rlabel alu0 278 105 278 105 1 a1b2_inv_1
rlabel alu1 247 152 247 152 6 vss
rlabel alu1 247 216 247 216 6 vdd
rlabel alu1 263 196 263 196 1 b1
rlabel alu1 255 188 255 188 1 b1
rlabel alu1 247 180 247 180 1 a2
rlabel alu1 255 176 255 176 1 a2
rlabel alu1 231 180 231 180 1 a2b1
rlabel alu0 252 200 252 200 1 a2b1_inv_0
rlabel alu0 239 183 239 183 1 a2b1_inv_0
rlabel alu1 164 117 164 117 1 a2b1
rlabel alu1 172 125 172 125 1 a2b1
rlabel alu1 245 113 245 113 1 a2b1
rlabel alu1 237 101 237 101 1 a2b1
rlabel alu0 227 105 227 105 1 a2b1_inv_1
rlabel alu0 242 132 242 132 1 a2b1_inv_1
rlabel alu1 53 145 53 145 2 vss
rlabel alu1 53 81 53 81 2 vdd
rlabel alu1 17 105 17 105 1 c04
rlabel ndifct1 17 133 17 133 1 c04
rlabel alu1 25 133 25 133 1 c04
rlabel alu1 33 133 33 133 1 c04
rlabel alu0 25 113 25 113 1 c04_inv_1
rlabel alu0 43 101 43 101 1 c04_inv_1
rlabel alu0 38 97 38 97 1 c04_inv_1
rlabel alu0 594 130 594 130 1 ha11
rlabel alu0 83 108 83 108 1 c04_inv_1
rlabel alu0 44 133 44 133 1 c04_inv_1
rlabel alu0 56 130 56 130 1 ha12
rlabel alu0 67 134 67 134 1 ha12
rlabel alu1 97 117 97 117 1 s04
rlabel alu1 89 93 89 93 1 s04
rlabel alu0 71 126 71 126 1 s04_inv_1
rlabel alu0 83 124 83 124 1 s04_inv_1
rlabel alu0 73 107 73 107 1 s04_inv_1
rlabel alu1 239 164 239 164 1 a2b1
rlabel alu1 100 152 100 152 6 vss
rlabel alu1 100 216 100 216 6 vdd
rlabel alu1 60 152 60 152 6 vss
rlabel alu1 60 216 60 216 6 vdd
rlabel alu1 116 196 116 196 1 b3
rlabel alu1 108 188 108 188 1 b3
rlabel alu1 100 180 100 180 1 a1
rlabel alu1 108 176 108 176 1 a1
rlabel alu1 84 180 84 180 1 a1b3
rlabel alu1 92 164 92 164 1 a1b3
rlabel alu0 105 200 105 200 1 a1b3_inv_0
rlabel alu0 92 183 92 183 1 a1b3_inv_0
rlabel alu0 108 164 108 164 1 a1b3_inv_0
rlabel alu1 65 113 65 113 1 a1b3
rlabel alu1 57 109 57 109 1 a1b3
rlabel alu1 49 109 49 109 1 a1b3
rlabel alu1 41 109 41 109 1 a1b3
rlabel alu1 33 109 33 109 1 a1b3
rlabel alu1 60 180 60 180 1 a2
rlabel alu1 68 176 68 176 1 a2
rlabel alu1 68 188 68 188 1 b2
rlabel alu1 76 196 76 196 1 b2
rlabel alu1 44 180 44 180 1 a2b2
rlabel alu0 65 200 65 200 1 a2b2_inv_0
rlabel alu0 52 183 52 183 1 a2b2_inv_0
rlabel alu0 68 164 68 164 1 a2b2_inv_0
rlabel alu1 52 164 52 164 1 a2b2
rlabel alu1 49 121 49 121 1 a2b2
rlabel alu1 41 117 41 117 1 a2b2
rlabel alu1 550 9 550 9 4 vss
rlabel alu1 550 73 550 73 4 vdd
rlabel alu1 514 49 514 49 1 c11
rlabel ndifct1 514 21 514 21 1 c11
rlabel alu1 522 21 522 21 1 c11
rlabel alu1 530 21 530 21 1 c11
rlabel alu0 535 57 535 57 1 c11_inv_2
rlabel alu0 540 53 540 53 1 c11_inv_2
rlabel alu0 522 41 522 41 1 c11_inv_2
rlabel alu0 580 46 580 46 1 c11_inv_2
rlabel alu1 594 37 594 37 1 res2
rlabel alu0 580 30 580 30 1 res2_inv
rlabel alu0 568 28 568 28 1 res2_inv
rlabel alu0 553 24 553 24 1 ha21
rlabel alu0 564 20 564 20 1 ha21
rlabel alu1 530 45 530 45 1 c01
rlabel alu1 538 45 538 45 1 c01
rlabel alu1 546 45 546 45 1 c01
rlabel alu1 562 41 562 41 1 c01
rlabel alu1 546 33 546 33 1 s02
rlabel alu0 541 21 541 21 1 c11_inv_2
rlabel alu0 570 47 570 47 1 res2_inv
rlabel alu1 586 61 586 61 1 res2
rlabel alu1 300 9 300 9 6 vss
rlabel alu1 300 73 300 73 6 vdd
rlabel alu1 344 9 344 9 6 vss
rlabel alu1 344 73 344 73 6 vdd
rlabel alu1 441 9 441 9 6 vss
rlabel alu1 441 73 441 73 6 vdd
rlabel alu1 292 37 292 37 1 c12
rlabel alu1 300 53 300 53 1 c12
rlabel alu1 308 37 308 37 1 c12_inv_2
rlabel alu1 300 33 300 33 1 c12_inv_2
rlabel alu1 340 29 340 29 1 c12_inv_2
rlabel alu0 320 57 320 57 1 fa_21_n1
rlabel alu0 348 62 348 62 1 fa_21_n1
rlabel alu0 336 20 336 20 1 fa_21_n3
rlabel alu0 356 21 356 21 1 fa_21_n3
rlabel alu1 389 53 389 53 1 s12
rlabel alu1 381 37 381 37 1 s12
rlabel alu1 389 21 389 21 1 s12
rlabel alu1 397 21 397 21 1 s12
rlabel alu1 316 41 316 41 1 s03
rlabel alu1 485 33 485 33 1 s03
rlabel polyct0 449 37 449 37 1 s03_inv_2
rlabel alu0 472 25 472 25 1 s03_inv_2
rlabel alu1 501 50 501 50 1 a3b0
rlabel alu1 364 41 364 41 1 a3b0
rlabel alu0 463 37 463 37 1 a3b0_inv_2
rlabel alu0 483 49 483 49 1 a3b0_inv_2
rlabel alu1 356 29 356 29 1 c02
rlabel alu1 429 41 429 41 1 c02
rlabel alu1 421 53 421 53 1 c02
rlabel alu0 411 49 411 49 1 c02_inv_2
rlabel alu0 426 22 426 22 1 c02_inv_2
rlabel alu0 462 49 462 49 1 s03_inv_2
rlabel alu0 493 36 493 36 1 a3b0_inv_2
rlabel alu1 143 216 143 216 6 vdd
rlabel alu1 143 152 143 152 6 vss
rlabel alu1 143 180 143 180 1 a3
rlabel alu0 454 164 454 164 1 a3b0_inv_0
rlabel alu1 151 188 151 188 1 b1
rlabel alu1 159 196 159 196 1 b1
rlabel alu1 127 180 127 180 1 a3b1
rlabel alu1 135 164 135 164 1 a3b1
rlabel alu0 135 183 135 183 1 a3b1_inv_0
rlabel alu1 80 9 80 9 6 vss
rlabel alu1 80 73 80 73 6 vdd
rlabel alu1 124 9 124 9 6 vss
rlabel alu1 124 73 124 73 6 vdd
rlabel alu1 221 9 221 9 6 vss
rlabel alu1 221 73 221 73 6 vdd
rlabel alu1 80 53 80 53 1 c13
rlabel alu1 72 37 72 37 1 c13
rlabel alu1 88 37 88 37 1 c13_inv_2
rlabel alu1 80 33 80 33 1 c13_inv_2
rlabel alu1 120 29 120 29 1 c13_inv_2
rlabel alu1 161 37 161 37 1 s13
rlabel alu1 169 53 169 53 1 s13
rlabel alu1 169 21 169 21 1 s13
rlabel alu1 177 21 177 21 1 s13
rlabel alu0 128 62 128 62 1 fa_22_n1
rlabel alu0 100 57 100 57 1 fa_22_n1
rlabel alu0 116 20 116 20 1 fa_22_n3
rlabel alu0 136 21 136 21 1 fa_22_n3
rlabel alu1 96 41 96 41 1 s04
rlabel alu1 265 33 265 33 1 s04
rlabel alu0 252 25 252 25 1 s04_inv_2
rlabel polyct0 229 37 229 37 1 s04_inv_2
rlabel alu0 242 49 242 49 1 s04_inv_2
rlabel alu1 144 41 144 41 1 c03
rlabel polyct1 281 45 281 45 1 c03
rlabel alu0 273 36 273 36 1 c03_inv_2
rlabel alu0 263 49 263 49 1 c03_inv_2
rlabel alu0 243 37 243 37 1 c03_inv_2
rlabel alu1 136 29 136 29 1 a3b1
rlabel alu1 128 37 128 37 1 a3b1
rlabel alu1 209 41 209 41 1 a3b1
rlabel alu1 201 53 201 53 1 a3b1
rlabel alu0 191 49 191 49 1 a3b1_inv_2
rlabel alu0 206 22 206 22 1 a3b1_inv_2
rlabel alu1 3 73 3 73 6 vdd
rlabel alu1 3 9 3 9 6 vss
rlabel alu1 -94 73 -94 73 6 vdd
rlabel alu1 -94 9 -94 9 6 vss
rlabel alu1 -138 73 -138 73 6 vdd
rlabel alu1 -138 9 -138 9 6 vss
rlabel alu1 -138 53 -138 53 1 c14
rlabel alu1 -146 37 -146 37 1 c14
rlabel alu1 -130 37 -130 37 1 c14_inv_2
rlabel alu1 -138 33 -138 33 1 c14_inv_2
rlabel alu1 -98 29 -98 29 1 c14_inv_2
rlabel alu0 -118 57 -118 57 1 fa_23_n1
rlabel alu0 -90 62 -90 62 1 fa_23_n1
rlabel alu0 -102 20 -102 20 1 fa_23_n3
rlabel alu0 -82 21 -82 21 1 fa_23_n3
rlabel alu1 -49 53 -49 53 1 s14
rlabel alu1 -57 37 -57 37 1 s14
rlabel alu1 -49 21 -49 21 1 s14
rlabel alu1 -41 21 -41 21 1 s14
rlabel alu1 -15 145 -15 145 8 vss
rlabel alu1 -15 81 -15 81 8 vdd
rlabel alu1 -57 81 -57 81 8 vdd
rlabel alu1 -57 145 -57 145 8 vss
rlabel alu1 -65 133 -65 133 1 a2b3
rlabel alu1 -73 117 -73 117 1 a2b3
rlabel alu0 -65 114 -65 114 1 a2b3_inv_1
rlabel alu0 -52 97 -52 97 1 a2b3_inv_1
rlabel alu1 -49 121 -49 121 1 a2
rlabel alu1 -57 117 -57 117 1 a2
rlabel alu1 -49 109 -49 109 1 b3
rlabel alu1 -41 101 -41 101 1 b3
rlabel alu1 -31 117 -31 117 1 a3b2
rlabel alu1 -23 133 -23 133 1 a3b2
rlabel alu0 -23 114 -23 114 1 a3b2_inv_1
rlabel alu0 -10 97 -10 97 1 a3b2_inv_1
rlabel alu1 -7 121 -7 121 1 a3
rlabel alu1 -15 117 -15 117 1 a3
rlabel alu1 -7 109 -7 109 1 b2
rlabel alu1 1 101 1 101 1 b2
rlabel alu0 -49 133 -49 133 1 a2b3_inv_1
rlabel alu0 -7 133 -7 133 1 a3b2_inv_1
rlabel alu1 -74 41 -74 41 1 a2b3
rlabel polyct1 63 45 63 45 1 a2b3
rlabel alu0 45 49 45 49 1 a2b3_inv_2
rlabel alu0 55 36 55 36 1 a2b3_inv_2
rlabel alu1 -122 41 -122 41 1 a3b2
rlabel alu1 47 33 47 33 1 a3b2
rlabel alu0 24 49 24 49 1 a3b2_inv_2
rlabel polyct0 11 37 11 37 1 a3b2_inv_2
rlabel alu0 34 25 34 25 1 a3b2_inv_2
rlabel alu1 -90 37 -90 37 1 c04
rlabel alu1 -82 29 -82 29 1 c04
rlabel alu1 -9 41 -9 41 1 c04
rlabel alu1 -17 53 -17 53 1 c04
rlabel alu0 -12 22 -12 22 1 c04_inv_2
rlabel alu0 -27 49 -27 49 1 c04_inv_2
rlabel alu1 493 -63 493 -63 2 vdd
rlabel alu1 493 1 493 1 2 vss
rlabel alu1 457 -39 457 -39 1 c21
rlabel ndifct1 457 -11 457 -11 1 c21
rlabel alu1 465 -11 465 -11 1 c21
rlabel alu1 473 -11 473 -11 1 c21
rlabel alu0 484 -11 484 -11 1 c21_inv_3
rlabel alu0 465 -31 465 -31 1 c21_inv_3
rlabel alu0 483 -43 483 -43 1 c21_inv_3
rlabel alu0 478 -47 478 -47 1 c21_inv_3
rlabel alu1 537 -27 537 -27 1 res3
rlabel alu1 529 -51 529 -51 1 res3
rlabel alu0 523 -36 523 -36 1 c21_inv_3
rlabel alu0 496 -14 496 -14 1 ha_31
rlabel alu0 507 -10 507 -10 1 ha_31
rlabel alu0 523 -20 523 -20 1 res3_inv
rlabel alu0 513 -37 513 -37 1 res3_inv
rlabel alu0 511 -18 511 -18 1 res3_inv
rlabel alu1 489 -23 489 -23 1 c11
rlabel alu1 481 -27 481 -27 1 c11
rlabel alu1 481 -35 481 -35 1 s12
rlabel alu1 489 -35 489 -35 1 s12
rlabel alu1 497 -35 497 -35 1 s12
rlabel alu1 505 -31 505 -31 1 s12
rlabel alu1 378 -63 378 -63 8 vdd
rlabel alu1 378 1 378 1 8 vss
rlabel alu1 281 -63 281 -63 8 vdd
rlabel alu1 281 1 281 1 8 vss
rlabel alu1 237 -63 237 -63 8 vdd
rlabel alu1 237 1 237 1 8 vss
rlabel alu0 273 -10 273 -10 1 fa_31_n3
rlabel alu0 293 -11 293 -11 1 fa_31_n3
rlabel alu0 257 -47 257 -47 1 fa_31_n1
rlabel alu0 285 -52 285 -52 1 fa_31_n1
rlabel alu1 318 -27 318 -27 1 res4
rlabel alu1 326 -43 326 -43 1 res4
rlabel alu1 326 -11 326 -11 1 res4
rlabel alu1 334 -11 334 -11 1 res4
rlabel polyct1 438 -35 438 -35 1 c21
rlabel via1 430 -43 430 -43 1 c21
rlabel via1 293 -43 293 -43 1 c21
rlabel alu1 301 -31 301 -31 1 c21
rlabel alu0 400 -27 400 -27 1 c21_inv_3_in
rlabel alu0 420 -39 420 -39 1 c21_inv_3_in
rlabel alu0 430 -26 430 -26 1 c21_inv_3_in
rlabel via1 301 -19 301 -19 1 c12
rlabel via1 293 -19 293 -19 1 c12
rlabel alu1 285 -27 285 -27 1 c12
rlabel alu1 366 -31 366 -31 1 c12
rlabel alu1 358 -43 358 -43 1 c12
rlabel alu0 363 -12 363 -12 1 c12_inv_3
rlabel alu0 348 -39 348 -39 1 c12_inv_3
rlabel via1 261 -27 261 -27 1 s13
rlabel alu1 253 -31 253 -31 1 s13
rlabel via1 414 -27 414 -27 1 s13
rlabel alu1 422 -23 422 -23 1 s13
rlabel polyct0 386 -27 386 -27 1 s13_inv_3
rlabel alu0 399 -39 399 -39 1 s13_inv_3
rlabel alu0 409 -15 409 -15 1 s13_inv_3
rlabel alu1 229 -27 229 -27 1 c22
rlabel alu1 277 -19 277 -19 1 c22_inv_3
rlabel alu1 245 -27 245 -27 1 c22_inv_3
rlabel alu1 237 -23 237 -23 1 c22_inv_3
rlabel alu1 237 -43 237 -43 1 c22
rlabel alu1 20 1 20 1 8 vss
rlabel alu1 20 -63 20 -63 8 vdd
rlabel alu1 64 1 64 1 8 vss
rlabel alu1 64 -63 64 -63 8 vdd
rlabel alu1 161 1 161 1 8 vss
rlabel alu1 161 -63 161 -63 8 vdd
rlabel alu1 12 -27 12 -27 1 c23
rlabel alu1 20 -43 20 -43 1 c23
rlabel alu1 20 -23 20 -23 1 c23_inv_3
rlabel alu1 28 -27 28 -27 1 c23_inv_3
rlabel alu1 60 -19 60 -19 1 c23_inv_3
rlabel alu0 56 -10 56 -10 1 fa_32_n3
rlabel alu0 76 -11 76 -11 1 fa_32_n3
rlabel alu0 40 -47 40 -47 1 fa_32_n1
rlabel alu0 68 -52 68 -52 1 fa_32_n1
rlabel alu1 101 -27 101 -27 1 res5
rlabel alu1 109 -43 109 -43 1 res5
rlabel alu1 109 -11 109 -11 1 res5
rlabel alu1 117 -11 117 -11 1 res5
rlabel polyct1 221 -35 221 -35 1 c22
rlabel via1 213 -43 213 -43 1 c22
rlabel via1 76 -43 76 -43 1 c22
rlabel alu1 84 -31 84 -31 1 c22
rlabel alu0 213 -26 213 -26 1 c22_inv_3_in
rlabel alu0 183 -27 183 -27 1 c22_inv_3_in
rlabel alu0 203 -39 203 -39 1 c22_inv_3_in
rlabel alu1 76 -19 76 -19 1 c13
rlabel via1 84 -19 84 -19 1 c13
rlabel alu1 68 -27 68 -27 1 c13
rlabel alu1 149 -31 149 -31 1 c13
rlabel alu1 141 -43 141 -43 1 c13
rlabel alu0 146 -12 146 -12 1 c13_inv_3
rlabel alu0 131 -39 131 -39 1 c13_inv_3
rlabel via1 44 -27 44 -27 1 s14
rlabel alu1 36 -31 36 -31 1 s14
rlabel via1 197 -27 197 -27 1 s14
rlabel alu1 205 -23 205 -23 1 s14
rlabel alu0 192 -15 192 -15 1 s14_inv_3
rlabel polyct0 169 -27 169 -27 1 s14_inv_3
rlabel alu0 182 -39 182 -39 1 s14_inv_3
rlabel alu1 -174 73 -174 73 6 vdd
rlabel alu1 -174 9 -174 9 6 vss
rlabel alu1 -190 37 -190 37 1 a3b3
rlabel alu1 -182 21 -182 21 1 a3b3
rlabel alu0 -169 57 -169 57 1 a3b3_inv_2
rlabel alu0 -182 40 -182 40 1 a3b3_inv_2
rlabel alu0 -166 21 -166 21 1 a3b3_inv_2
rlabel alu1 -174 37 -174 37 1 a3
rlabel alu1 -166 33 -166 33 1 a3
rlabel alu1 -166 45 -166 45 1 b3
rlabel alu1 -158 53 -158 53 1 b3
rlabel alu1 -59 -63 -59 -63 8 vdd
rlabel alu1 -59 1 -59 1 8 vss
rlabel alu1 -156 -63 -156 -63 8 vdd
rlabel alu1 -156 1 -156 1 8 vss
rlabel alu1 -200 -63 -200 -63 8 vdd
rlabel alu1 -200 1 -200 1 8 vss
rlabel alu1 -208 -27 -208 -27 1 res7
rlabel alu1 -200 -43 -200 -43 1 res7
rlabel alu1 -200 -23 -200 -23 1 res7_inv
rlabel alu1 -192 -27 -192 -27 1 res7_inv
rlabel alu1 -160 -19 -160 -19 1 res7_inv
rlabel alu0 -164 -10 -164 -10 1 fa_33_n3
rlabel alu0 -144 -11 -144 -11 1 fa_33_n3
rlabel alu0 -180 -47 -180 -47 1 fa_33_n1
rlabel alu0 -152 -52 -152 -52 1 fa_33_n1
rlabel alu1 -111 -43 -111 -43 1 res6
rlabel alu1 -119 -27 -119 -27 1 res6
rlabel alu1 -111 -11 -111 -11 1 res6
rlabel alu1 -103 -11 -103 -11 1 res6
rlabel polyct1 1 -35 1 -35 1 c23
rlabel via1 -7 -43 -7 -43 1 c23
rlabel via1 -144 -43 -144 -43 1 c23
rlabel alu1 -136 -31 -136 -31 1 c23
rlabel alu0 -7 -26 -7 -26 1 c23_inv_3_in
rlabel alu0 -17 -39 -17 -39 1 c23_inv_3_in
rlabel alu0 -37 -27 -37 -27 1 c23_inv_3_in
rlabel via1 -136 -19 -136 -19 1 c14
rlabel alu1 -144 -19 -144 -19 1 c14
rlabel alu1 -152 -27 -152 -27 1 c14
rlabel alu1 -71 -31 -71 -31 1 c14
rlabel alu1 -79 -43 -79 -43 1 c14
rlabel alu0 -74 -12 -74 -12 1 c14_inv_3
rlabel alu0 -89 -39 -89 -39 1 c14_inv_3
rlabel alu1 -184 -31 -184 -31 1 a3b3
rlabel via1 -176 -27 -176 -27 1 a3b3
rlabel via1 -23 -27 -23 -27 1 a3b3
rlabel alu1 -15 -23 -15 -23 1 a3b3
rlabel alu0 -28 -15 -28 -15 1 a3b3_inv_3
rlabel polyct0 -51 -27 -51 -27 1 a3b3_inv_3
rlabel alu0 -38 -39 -38 -39 1 a3b3_inv_3
<< end >>
